*cla_adder
.include TSMC_180nm.txt
.param LAMBDA = 0.09u
.param SUPPLY = 1.8v
.param W = {20*LAMBDA}
.param WIDTH_N = {W}
.param WIDTH_P = {2*W} 
.global gnd Vdd

VDD Vdd gnd DC 'SUPPLY'

Va0 x gnd PULSE(0 1.8 0ns 10ps 10ps 5ns 10ns)

.subckt inverter ip op vdd gnd S=1
.param w_p = {2*W}
.param w_n = {W}

Minv1 op ip vdd vdd CMOSP W={S*w_p} L={2*LAMBDA} 
+ AS={S*5*w_p*LAMBDA} PS={10*LAMBDA+S*2*w_p} 
+ AD={S*5*w_p*LAMBDA} PD={10*LAMBDA+S*2*w_p}

Minv2 op ip gnd gnd CMOSN W={S*w_n} L={2*LAMBDA} 
+ AS={S*5*w_n*LAMBDA} PS={10*LAMBDA+S*2*w_n} 
+ AD={S*5*w_n*LAMBDA} PD={10*LAMBDA+S*2*w_n}
.ends inverter

X1 x y vdd gnd inverter

.tran 1ps 20ns

.measure tran tpcq_inv
+TRIG v(x) VAL=0.9 FALL=1
+TARG v(y) VAL=0.9 RISE=1

.control
run
set color0 = white
set xbrushwidth = 3
set hcopypscolor=1
set curplottitle = "raviSahu2024102024_CLAADDER"
plot v(y) 4+v(x)
hardcopy inverter_plot.ps v(y) 4+v(x)
.endc