magic
tech scmos
timestamp 1764667915
<< error_p >>
rect 0 1 1 3
rect 0 0 3 1
<< nwell >>
rect -74 -654 -42 161
rect 22 69 54 136
rect 280 135 368 167
rect 22 21 76 69
rect 22 -63 54 21
rect 215 -22 247 15
rect 361 6 392 11
rect 361 -26 393 6
rect 22 -111 76 -63
rect 215 -98 247 -28
rect 498 -31 530 -7
rect 361 -97 393 -52
rect 498 -79 552 -31
rect 22 -198 54 -111
rect 22 -246 76 -198
rect 215 -215 247 -104
rect 498 -121 530 -79
rect 361 -202 393 -149
rect 498 -169 552 -121
rect 498 -210 530 -169
rect 22 -330 54 -246
rect 22 -378 76 -330
rect 22 -464 54 -378
rect 215 -381 247 -221
rect 498 -258 552 -210
rect 361 -352 394 -291
rect 498 -298 530 -258
rect 498 -346 552 -298
rect 498 -387 530 -346
rect 22 -512 76 -464
rect 22 -536 54 -512
rect 215 -604 247 -387
rect 498 -435 552 -387
rect 498 -459 530 -435
rect 628 -472 660 21
rect 361 -566 394 -497
<< ntransistor >>
rect -30 148 -20 150
rect -30 132 -20 134
rect -30 124 -20 126
rect 95 123 105 125
rect 291 113 293 123
rect 307 113 309 123
rect 315 113 317 123
rect 331 113 333 123
rect 339 113 341 123
rect 355 113 357 123
rect -30 108 -20 110
rect 87 106 107 108
rect -30 100 -20 102
rect 87 98 107 100
rect -30 84 -20 86
rect 90 80 100 82
rect -30 67 -20 69
rect 85 56 105 58
rect -30 51 -20 53
rect 85 48 105 50
rect -30 43 -20 45
rect 85 40 105 42
rect 85 32 105 34
rect -30 27 -20 29
rect -30 19 -20 21
rect 90 8 100 10
rect 672 8 682 10
rect -30 3 -20 5
rect 257 -3 277 -1
rect 95 -9 105 -7
rect -30 -13 -20 -11
rect 401 -7 421 -5
rect 257 -11 277 -9
rect 672 -8 682 -6
rect 401 -15 421 -13
rect -30 -29 -20 -27
rect 672 -16 682 -14
rect 566 -20 576 -18
rect 87 -26 107 -24
rect 87 -34 107 -32
rect -30 -37 -20 -35
rect 672 -32 682 -30
rect -30 -53 -20 -51
rect 672 -40 682 -38
rect 561 -44 581 -42
rect 257 -46 287 -44
rect 90 -52 100 -50
rect 561 -52 581 -50
rect 257 -54 287 -52
rect -30 -61 -20 -59
rect 257 -62 287 -60
rect 672 -56 682 -54
rect 561 -60 581 -58
rect 403 -70 433 -68
rect 561 -68 581 -66
rect -30 -77 -20 -75
rect 85 -76 105 -74
rect 257 -79 277 -77
rect 672 -73 682 -71
rect 403 -78 433 -76
rect 85 -84 105 -82
rect -30 -94 -20 -92
rect 257 -87 277 -85
rect 403 -86 433 -84
rect 85 -92 105 -90
rect 672 -89 682 -87
rect 566 -92 576 -90
rect 672 -97 682 -95
rect 85 -100 105 -98
rect -30 -110 -20 -108
rect 566 -110 576 -108
rect 672 -113 682 -111
rect -30 -118 -20 -116
rect 90 -124 100 -122
rect 256 -122 296 -120
rect 672 -121 682 -119
rect 256 -130 296 -128
rect -30 -134 -20 -132
rect -30 -142 -20 -140
rect 561 -134 581 -132
rect 256 -138 296 -136
rect 95 -144 105 -142
rect 672 -137 682 -135
rect 561 -142 581 -140
rect 256 -146 296 -144
rect 561 -150 581 -148
rect -30 -158 -20 -156
rect 87 -161 107 -159
rect 672 -154 682 -152
rect 561 -158 581 -156
rect 256 -163 286 -161
rect 87 -169 107 -167
rect -30 -175 -20 -173
rect 402 -167 432 -165
rect 256 -171 286 -169
rect 672 -170 682 -168
rect 402 -175 432 -173
rect 256 -179 286 -177
rect 402 -183 432 -181
rect 672 -178 682 -176
rect 566 -182 576 -180
rect 90 -187 100 -185
rect -30 -191 -20 -189
rect -30 -199 -20 -197
rect 402 -191 432 -189
rect 256 -196 276 -194
rect 672 -194 682 -192
rect 566 -199 576 -197
rect 256 -204 276 -202
rect 672 -202 682 -200
rect 85 -211 105 -209
rect -30 -215 -20 -213
rect 85 -219 105 -217
rect -30 -223 -20 -221
rect 672 -218 682 -216
rect 561 -223 581 -221
rect 85 -227 105 -225
rect 561 -231 581 -229
rect 85 -235 105 -233
rect -30 -239 -20 -237
rect 256 -239 306 -237
rect 672 -235 682 -233
rect 561 -239 581 -237
rect 256 -247 306 -245
rect -30 -256 -20 -254
rect 561 -247 581 -245
rect 672 -251 682 -249
rect 256 -255 306 -253
rect 90 -259 100 -257
rect 672 -259 682 -257
rect 256 -263 306 -261
rect -30 -272 -20 -270
rect 256 -271 306 -269
rect 95 -276 105 -274
rect 566 -271 576 -269
rect 672 -275 682 -273
rect -30 -280 -20 -278
rect -30 -296 -20 -294
rect 256 -288 296 -286
rect 672 -283 682 -281
rect 566 -287 576 -285
rect 87 -293 107 -291
rect 256 -296 296 -294
rect 87 -301 107 -299
rect -30 -304 -20 -302
rect 672 -299 682 -297
rect 256 -304 296 -302
rect -30 -320 -20 -318
rect 402 -309 442 -307
rect 256 -312 296 -310
rect 90 -319 100 -317
rect 561 -311 581 -309
rect 402 -317 442 -315
rect 672 -316 682 -314
rect 561 -319 581 -317
rect 402 -325 442 -323
rect 256 -329 286 -327
rect -30 -336 -20 -334
rect 561 -327 581 -325
rect 402 -333 442 -331
rect 256 -337 286 -335
rect 85 -343 105 -341
rect 672 -332 682 -330
rect 561 -335 581 -333
rect 402 -341 442 -339
rect 672 -340 682 -338
rect 256 -345 286 -343
rect -30 -352 -20 -350
rect 85 -351 105 -349
rect -30 -360 -20 -358
rect 85 -359 105 -357
rect 672 -356 682 -354
rect 566 -359 576 -357
rect 256 -362 276 -360
rect 85 -367 105 -365
rect 672 -364 682 -362
rect 256 -370 276 -368
rect -30 -376 -20 -374
rect 566 -376 576 -374
rect 672 -380 682 -378
rect -30 -384 -20 -382
rect 90 -391 100 -389
rect 672 -397 682 -395
rect -30 -400 -20 -398
rect 561 -400 581 -398
rect 256 -405 316 -403
rect 95 -410 105 -408
rect 561 -408 581 -406
rect 256 -413 316 -411
rect -30 -417 -20 -415
rect 672 -413 682 -411
rect 561 -416 581 -414
rect 256 -421 316 -419
rect 87 -427 107 -425
rect -30 -433 -20 -431
rect 672 -421 682 -419
rect 561 -424 581 -422
rect 256 -429 316 -427
rect 87 -435 107 -433
rect -30 -441 -20 -439
rect 256 -437 316 -435
rect 672 -437 682 -435
rect 256 -445 316 -443
rect 672 -445 682 -443
rect 566 -448 576 -446
rect 90 -453 100 -451
rect -30 -457 -20 -455
rect -30 -465 -20 -463
rect 256 -462 306 -460
rect 672 -461 682 -459
rect 256 -470 306 -468
rect 85 -477 105 -475
rect -30 -481 -20 -479
rect 256 -478 306 -476
rect 85 -485 105 -483
rect 256 -486 306 -484
rect 85 -493 105 -491
rect -30 -498 -20 -496
rect 256 -494 306 -492
rect 85 -501 105 -499
rect -30 -514 -20 -512
rect 256 -511 296 -509
rect -30 -522 -20 -520
rect 405 -515 465 -513
rect 256 -519 296 -517
rect 90 -525 100 -523
rect 405 -523 465 -521
rect 256 -527 296 -525
rect -30 -538 -20 -536
rect 405 -531 465 -529
rect 256 -535 296 -533
rect 405 -539 465 -537
rect -30 -546 -20 -544
rect 405 -547 465 -545
rect 256 -552 286 -550
rect -30 -562 -20 -560
rect 405 -555 465 -553
rect 256 -560 286 -558
rect 256 -568 286 -566
rect -30 -579 -20 -577
rect 256 -585 276 -583
rect -30 -595 -20 -593
rect 256 -593 276 -591
rect -30 -603 -20 -601
rect -30 -619 -20 -617
rect -30 -627 -20 -625
rect -30 -643 -20 -641
<< ptransistor >>
rect -68 148 -48 150
rect 291 141 293 161
rect 315 141 317 161
rect 331 141 333 161
rect 347 141 349 161
rect 355 141 357 161
rect -68 124 -48 126
rect 28 123 48 125
rect -68 108 -48 110
rect 28 106 48 108
rect 28 98 48 100
rect -68 92 -48 94
rect -68 84 -48 86
rect 28 80 48 82
rect -68 67 -48 69
rect 29 56 69 58
rect 29 48 69 50
rect -68 43 -48 45
rect 29 40 69 42
rect 29 32 69 34
rect -68 27 -48 29
rect -68 11 -48 13
rect 28 8 48 10
rect 634 8 654 10
rect -68 3 -48 5
rect 221 -3 241 -1
rect 28 -9 48 -7
rect -68 -13 -48 -11
rect 367 -7 387 -5
rect 221 -11 241 -9
rect 367 -15 387 -13
rect 634 -16 654 -14
rect 504 -20 524 -18
rect 28 -26 48 -24
rect 28 -34 48 -32
rect -68 -37 -48 -35
rect 634 -32 654 -30
rect -68 -53 -48 -51
rect 505 -44 545 -42
rect 221 -46 241 -44
rect 28 -52 48 -50
rect 634 -48 654 -46
rect 505 -52 545 -50
rect 221 -54 241 -52
rect 221 -62 241 -60
rect 634 -56 654 -54
rect 505 -60 545 -58
rect -68 -69 -48 -67
rect 367 -70 387 -68
rect 505 -68 545 -66
rect -68 -77 -48 -75
rect 29 -76 69 -74
rect 221 -79 241 -77
rect 634 -73 654 -71
rect 367 -78 387 -76
rect 29 -84 69 -82
rect -68 -94 -48 -92
rect 221 -87 241 -85
rect 367 -86 387 -84
rect 29 -92 69 -90
rect 504 -92 524 -90
rect 634 -97 654 -95
rect 29 -100 69 -98
rect 504 -110 524 -108
rect 634 -113 654 -111
rect -68 -118 -48 -116
rect 28 -124 48 -122
rect 221 -122 241 -120
rect 221 -130 241 -128
rect -68 -134 -48 -132
rect 634 -129 654 -127
rect 505 -134 545 -132
rect 221 -138 241 -136
rect 28 -144 48 -142
rect -68 -150 -48 -148
rect 634 -137 654 -135
rect 505 -142 545 -140
rect 221 -146 241 -144
rect 505 -150 545 -148
rect -68 -158 -48 -156
rect 28 -161 48 -159
rect 634 -154 654 -152
rect 505 -158 545 -156
rect 221 -163 241 -161
rect 28 -169 48 -167
rect -68 -175 -48 -173
rect 367 -167 387 -165
rect 221 -171 241 -169
rect 367 -175 387 -173
rect 221 -179 241 -177
rect 367 -183 387 -181
rect 634 -178 654 -176
rect 504 -182 524 -180
rect 28 -187 48 -185
rect -68 -199 -48 -197
rect 367 -191 387 -189
rect 221 -196 241 -194
rect 634 -194 654 -192
rect 504 -199 524 -197
rect 221 -204 241 -202
rect 29 -211 69 -209
rect -68 -215 -48 -213
rect 634 -210 654 -208
rect 29 -219 69 -217
rect 634 -218 654 -216
rect 505 -223 545 -221
rect 29 -227 69 -225
rect -68 -231 -48 -229
rect 505 -231 545 -229
rect 29 -235 69 -233
rect -68 -239 -48 -237
rect 221 -239 241 -237
rect 634 -235 654 -233
rect 505 -239 545 -237
rect 221 -247 241 -245
rect -68 -256 -48 -254
rect 505 -247 545 -245
rect 221 -255 241 -253
rect 28 -259 48 -257
rect 634 -259 654 -257
rect 221 -263 241 -261
rect 221 -271 241 -269
rect 28 -276 48 -274
rect 504 -271 524 -269
rect 634 -275 654 -273
rect -68 -280 -48 -278
rect -68 -296 -48 -294
rect 221 -288 241 -286
rect 504 -287 524 -285
rect 28 -293 48 -291
rect 634 -291 654 -289
rect 221 -296 241 -294
rect 28 -301 48 -299
rect 634 -299 654 -297
rect 221 -304 241 -302
rect -68 -312 -48 -310
rect -68 -320 -48 -318
rect 368 -309 388 -307
rect 221 -312 241 -310
rect 28 -319 48 -317
rect 505 -311 545 -309
rect 368 -317 388 -315
rect 634 -316 654 -314
rect 505 -319 545 -317
rect 368 -325 388 -323
rect 221 -329 241 -327
rect -68 -336 -48 -334
rect 505 -327 545 -325
rect 368 -333 388 -331
rect 221 -337 241 -335
rect 29 -343 69 -341
rect 505 -335 545 -333
rect 368 -341 388 -339
rect 634 -340 654 -338
rect 221 -345 241 -343
rect 29 -351 69 -349
rect -68 -360 -48 -358
rect 29 -359 69 -357
rect 634 -356 654 -354
rect 504 -359 524 -357
rect 221 -362 241 -360
rect 29 -367 69 -365
rect 221 -370 241 -368
rect -68 -376 -48 -374
rect 634 -372 654 -370
rect 504 -376 524 -374
rect 634 -380 654 -378
rect -68 -392 -48 -390
rect 28 -391 48 -389
rect 634 -397 654 -395
rect -68 -400 -48 -398
rect 505 -400 545 -398
rect 221 -405 241 -403
rect 28 -410 48 -408
rect 505 -408 545 -406
rect 221 -413 241 -411
rect -68 -417 -48 -415
rect 505 -416 545 -414
rect 221 -421 241 -419
rect 28 -427 48 -425
rect 634 -421 654 -419
rect 505 -424 545 -422
rect 221 -429 241 -427
rect 28 -435 48 -433
rect -68 -441 -48 -439
rect 221 -437 241 -435
rect 634 -437 654 -435
rect 221 -445 241 -443
rect 504 -448 524 -446
rect 28 -453 48 -451
rect -68 -457 -48 -455
rect 634 -453 654 -451
rect 221 -462 241 -460
rect 634 -461 654 -459
rect -68 -473 -48 -471
rect 221 -470 241 -468
rect 29 -477 69 -475
rect -68 -481 -48 -479
rect 221 -478 241 -476
rect 29 -485 69 -483
rect 221 -486 241 -484
rect 29 -493 69 -491
rect -68 -498 -48 -496
rect 221 -494 241 -492
rect 29 -501 69 -499
rect 221 -511 241 -509
rect -68 -522 -48 -520
rect 368 -515 388 -513
rect 221 -519 241 -517
rect 28 -525 48 -523
rect 368 -523 388 -521
rect 221 -527 241 -525
rect -68 -538 -48 -536
rect 368 -531 388 -529
rect 221 -535 241 -533
rect 368 -539 388 -537
rect -68 -554 -48 -552
rect 368 -547 388 -545
rect 221 -552 241 -550
rect -68 -562 -48 -560
rect 368 -555 388 -553
rect 221 -560 241 -558
rect 221 -568 241 -566
rect -68 -579 -48 -577
rect 221 -585 241 -583
rect 221 -593 241 -591
rect -68 -603 -48 -601
rect -68 -619 -48 -617
rect -68 -635 -48 -633
rect -68 -643 -48 -641
<< ndiffusion >>
rect -26 151 -20 155
rect -30 150 -20 151
rect -30 147 -20 148
rect -30 143 -24 147
rect -26 135 -20 139
rect -30 134 -20 135
rect -30 126 -20 132
rect 99 126 105 130
rect 95 125 105 126
rect -30 123 -20 124
rect -30 119 -24 123
rect 95 122 105 123
rect 95 118 101 122
rect 290 119 291 123
rect -30 111 -24 115
rect 286 113 291 119
rect 293 117 298 123
rect 293 113 294 117
rect 306 119 307 123
rect 302 113 307 119
rect 309 113 315 123
rect 317 117 322 123
rect 317 113 318 117
rect 326 117 331 123
rect 330 113 331 117
rect 333 113 339 123
rect 341 119 342 123
rect 341 113 346 119
rect 354 119 355 123
rect 350 113 355 119
rect 357 117 362 123
rect 357 113 358 117
rect -30 110 -20 111
rect -30 102 -20 108
rect 91 109 107 113
rect 87 108 107 109
rect -30 99 -20 100
rect -26 95 -20 99
rect 87 100 107 106
rect 87 97 107 98
rect 87 93 103 97
rect -26 87 -20 91
rect -30 86 -20 87
rect -30 83 -20 84
rect -30 79 -24 83
rect 90 83 96 87
rect 90 82 100 83
rect 90 79 100 80
rect 94 75 100 79
rect -26 70 -20 74
rect -30 69 -20 70
rect -30 66 -20 67
rect -30 62 -24 66
rect 89 59 105 63
rect 85 58 105 59
rect -26 54 -20 58
rect -30 53 -20 54
rect -30 45 -20 51
rect 85 50 105 56
rect -30 42 -20 43
rect -30 38 -24 42
rect 85 47 105 48
rect 85 43 101 47
rect 85 42 105 43
rect -30 30 -24 34
rect 85 34 105 40
rect -30 29 -20 30
rect -30 21 -20 27
rect 85 31 105 32
rect 89 27 105 31
rect -30 18 -20 19
rect -26 14 -20 18
rect -26 6 -20 10
rect 94 11 100 15
rect 90 10 100 11
rect 676 11 682 15
rect 672 10 682 11
rect -30 5 -20 6
rect 90 7 100 8
rect 90 3 96 7
rect -30 2 -20 3
rect -30 -2 -24 2
rect -26 -10 -20 -6
rect 99 -6 105 -2
rect 257 0 273 4
rect 672 7 682 8
rect 672 3 678 7
rect 257 -1 277 0
rect 95 -7 105 -6
rect -30 -11 -20 -10
rect -30 -14 -20 -13
rect 95 -10 105 -9
rect 95 -14 101 -10
rect 257 -9 277 -3
rect 401 -4 417 0
rect 401 -5 421 -4
rect 676 -5 682 -1
rect 672 -6 682 -5
rect -30 -18 -24 -14
rect 257 -12 277 -11
rect 261 -16 277 -12
rect 401 -13 421 -7
rect -26 -26 -20 -22
rect -30 -27 -20 -26
rect -30 -35 -20 -29
rect 91 -23 107 -19
rect 401 -16 421 -15
rect 405 -20 421 -16
rect 566 -17 572 -13
rect 672 -14 682 -8
rect 566 -18 576 -17
rect 87 -24 107 -23
rect 566 -21 576 -20
rect 672 -17 682 -16
rect 672 -21 678 -17
rect 570 -25 576 -21
rect 87 -32 107 -26
rect -30 -38 -20 -37
rect -30 -42 -24 -38
rect 87 -35 107 -34
rect 672 -29 678 -25
rect 672 -30 682 -29
rect 87 -39 103 -35
rect -30 -50 -24 -46
rect -30 -51 -20 -50
rect -30 -59 -20 -53
rect 90 -49 96 -45
rect 257 -43 283 -39
rect 565 -41 581 -37
rect 672 -38 682 -32
rect 672 -41 682 -40
rect 561 -42 581 -41
rect 257 -44 287 -43
rect 90 -50 100 -49
rect 90 -53 100 -52
rect 94 -57 100 -53
rect 257 -52 287 -46
rect 561 -50 581 -44
rect 676 -45 682 -41
rect -30 -62 -20 -61
rect -26 -66 -20 -62
rect 257 -60 287 -54
rect 561 -53 581 -52
rect 561 -57 577 -53
rect 676 -53 682 -49
rect 672 -54 682 -53
rect 561 -58 581 -57
rect 257 -63 287 -62
rect 261 -67 287 -63
rect -26 -74 -20 -70
rect 89 -73 105 -69
rect 403 -67 429 -63
rect 403 -68 433 -67
rect 561 -66 581 -60
rect 672 -57 682 -56
rect 672 -61 678 -57
rect 85 -74 105 -73
rect -30 -75 -20 -74
rect -30 -78 -20 -77
rect -30 -82 -24 -78
rect 85 -82 105 -76
rect 257 -76 273 -72
rect 257 -77 277 -76
rect 403 -76 433 -70
rect 561 -69 581 -68
rect 565 -73 581 -69
rect 676 -70 682 -66
rect 672 -71 682 -70
rect 672 -74 682 -73
rect 672 -78 678 -74
rect -26 -91 -20 -87
rect -30 -92 -20 -91
rect 85 -85 105 -84
rect 85 -89 101 -85
rect 257 -85 277 -79
rect 403 -84 433 -78
rect 85 -90 105 -89
rect 257 -88 277 -87
rect 261 -92 277 -88
rect 403 -87 433 -86
rect 407 -91 433 -87
rect -30 -95 -20 -94
rect -30 -99 -24 -95
rect 85 -98 105 -92
rect 570 -89 576 -85
rect 676 -86 682 -82
rect 672 -87 682 -86
rect 566 -90 576 -89
rect 566 -93 576 -92
rect 566 -97 572 -93
rect 672 -95 682 -89
rect -26 -107 -20 -103
rect 85 -101 105 -100
rect 89 -105 105 -101
rect 672 -98 682 -97
rect 672 -102 678 -98
rect -30 -108 -20 -107
rect -30 -116 -20 -110
rect 566 -107 572 -103
rect 566 -108 576 -107
rect 566 -111 576 -110
rect 570 -115 576 -111
rect 672 -110 678 -106
rect 672 -111 682 -110
rect -30 -119 -20 -118
rect -30 -123 -24 -119
rect 94 -121 100 -117
rect 90 -122 100 -121
rect 256 -119 292 -115
rect 256 -120 296 -119
rect -30 -131 -24 -127
rect 90 -125 100 -124
rect 90 -129 96 -125
rect 256 -128 296 -122
rect 672 -119 682 -113
rect 672 -122 682 -121
rect 676 -126 682 -122
rect -30 -132 -20 -131
rect -30 -140 -20 -134
rect 99 -141 105 -137
rect 256 -136 296 -130
rect 565 -131 581 -127
rect 561 -132 581 -131
rect 95 -142 105 -141
rect -30 -143 -20 -142
rect -26 -147 -20 -143
rect 95 -145 105 -144
rect 95 -149 101 -145
rect 256 -144 296 -138
rect 561 -140 581 -134
rect 676 -134 682 -130
rect 672 -135 682 -134
rect 256 -147 296 -146
rect 260 -151 296 -147
rect 561 -143 581 -142
rect 672 -138 682 -137
rect 672 -142 678 -138
rect 561 -147 577 -143
rect 561 -148 581 -147
rect -26 -155 -20 -151
rect -30 -156 -20 -155
rect -30 -159 -20 -158
rect -30 -163 -24 -159
rect 91 -158 107 -154
rect 87 -159 107 -158
rect -26 -172 -20 -168
rect 87 -167 107 -161
rect 256 -160 282 -156
rect 561 -156 581 -150
rect 676 -151 682 -147
rect 672 -152 682 -151
rect 256 -161 286 -160
rect -30 -173 -20 -172
rect 87 -170 107 -169
rect 87 -174 103 -170
rect 256 -169 286 -163
rect 402 -164 428 -160
rect 561 -159 581 -158
rect 672 -155 682 -154
rect 672 -159 678 -155
rect 565 -163 581 -159
rect 402 -165 432 -164
rect 676 -167 682 -163
rect -30 -176 -20 -175
rect -30 -180 -24 -176
rect 256 -177 286 -171
rect 402 -173 432 -167
rect 672 -168 682 -167
rect -26 -188 -20 -184
rect 90 -184 96 -180
rect 256 -180 286 -179
rect 260 -184 286 -180
rect 402 -181 432 -175
rect 570 -179 576 -175
rect 672 -176 682 -170
rect 566 -180 576 -179
rect 90 -185 100 -184
rect -30 -189 -20 -188
rect -30 -197 -20 -191
rect 90 -188 100 -187
rect 94 -192 100 -188
rect -30 -200 -20 -199
rect 256 -193 272 -189
rect 402 -189 432 -183
rect 566 -183 576 -182
rect 672 -179 682 -178
rect 672 -183 678 -179
rect 566 -187 572 -183
rect 256 -194 276 -193
rect 402 -192 432 -191
rect 406 -196 432 -192
rect -30 -204 -24 -200
rect -30 -212 -24 -208
rect 89 -208 105 -204
rect 256 -202 276 -196
rect 566 -196 572 -192
rect 672 -191 678 -187
rect 672 -192 682 -191
rect 566 -197 576 -196
rect 566 -200 576 -199
rect 570 -204 576 -200
rect 672 -200 682 -194
rect 672 -203 682 -202
rect 85 -209 105 -208
rect -30 -213 -20 -212
rect -30 -221 -20 -215
rect 85 -217 105 -211
rect 256 -205 276 -204
rect 260 -209 276 -205
rect 676 -207 682 -203
rect -30 -224 -20 -223
rect -26 -228 -20 -224
rect 85 -220 105 -219
rect 85 -224 101 -220
rect 565 -220 581 -216
rect 676 -215 682 -211
rect 672 -216 682 -215
rect 561 -221 581 -220
rect 85 -225 105 -224
rect -26 -236 -20 -232
rect 85 -233 105 -227
rect 561 -229 581 -223
rect 672 -219 682 -218
rect 672 -223 678 -219
rect -30 -237 -20 -236
rect -30 -240 -20 -239
rect 85 -236 105 -235
rect 89 -240 105 -236
rect 256 -236 302 -232
rect 256 -237 306 -236
rect -30 -244 -24 -240
rect 256 -245 306 -239
rect 561 -232 581 -231
rect 561 -236 577 -232
rect 676 -232 682 -228
rect 672 -233 682 -232
rect 561 -237 581 -236
rect -26 -253 -20 -249
rect -30 -254 -20 -253
rect -30 -257 -20 -256
rect -30 -261 -24 -257
rect 94 -256 100 -252
rect 256 -253 306 -247
rect 561 -245 581 -239
rect 672 -236 682 -235
rect 672 -240 678 -236
rect 561 -248 581 -247
rect 676 -248 682 -244
rect 565 -252 581 -248
rect 672 -249 682 -248
rect 90 -257 100 -256
rect 90 -260 100 -259
rect 90 -264 96 -260
rect 256 -261 306 -255
rect 672 -257 682 -251
rect -26 -269 -20 -265
rect -30 -270 -20 -269
rect -30 -278 -20 -272
rect 99 -273 105 -269
rect 256 -269 306 -263
rect 672 -260 682 -259
rect 672 -264 678 -260
rect 95 -274 105 -273
rect 256 -272 306 -271
rect 570 -268 576 -264
rect 566 -269 576 -268
rect 260 -276 306 -272
rect 566 -272 576 -271
rect 566 -276 572 -272
rect 672 -272 678 -268
rect 672 -273 682 -272
rect -30 -281 -20 -280
rect 95 -277 105 -276
rect 95 -281 101 -277
rect -30 -285 -24 -281
rect -30 -293 -24 -289
rect -30 -294 -20 -293
rect -30 -302 -20 -296
rect 91 -290 107 -286
rect 256 -285 292 -281
rect 256 -286 296 -285
rect 566 -284 572 -280
rect 672 -281 682 -275
rect 672 -284 682 -283
rect 566 -285 576 -284
rect 87 -291 107 -290
rect 87 -299 107 -293
rect 256 -294 296 -288
rect 566 -288 576 -287
rect 676 -288 682 -284
rect 570 -292 576 -288
rect -30 -305 -20 -304
rect -26 -309 -20 -305
rect 87 -302 107 -301
rect 87 -306 103 -302
rect 256 -302 296 -296
rect 676 -296 682 -292
rect 672 -297 682 -296
rect -26 -317 -20 -313
rect -30 -318 -20 -317
rect 90 -316 96 -312
rect 256 -310 296 -304
rect 402 -306 438 -302
rect 672 -300 682 -299
rect 672 -304 678 -300
rect 402 -307 442 -306
rect 565 -308 581 -304
rect 561 -309 581 -308
rect 90 -317 100 -316
rect 256 -313 296 -312
rect 260 -317 296 -313
rect 402 -315 442 -309
rect 561 -317 581 -311
rect 676 -313 682 -309
rect 672 -314 682 -313
rect -30 -321 -20 -320
rect -30 -325 -24 -321
rect 90 -320 100 -319
rect 94 -324 100 -320
rect -26 -333 -20 -329
rect 256 -326 282 -322
rect 402 -323 442 -317
rect 256 -327 286 -326
rect -30 -334 -20 -333
rect -30 -337 -20 -336
rect -30 -341 -24 -337
rect 89 -340 105 -336
rect 256 -335 286 -329
rect 402 -331 442 -325
rect 561 -320 581 -319
rect 561 -324 577 -320
rect 672 -317 682 -316
rect 672 -321 678 -317
rect 561 -325 581 -324
rect 85 -341 105 -340
rect -26 -349 -20 -345
rect 85 -349 105 -343
rect 256 -343 286 -337
rect 402 -339 442 -333
rect 561 -333 581 -327
rect 676 -329 682 -325
rect 672 -330 682 -329
rect 561 -336 581 -335
rect 565 -340 581 -336
rect 672 -338 682 -332
rect -30 -350 -20 -349
rect -30 -358 -20 -352
rect 85 -352 105 -351
rect 256 -346 286 -345
rect 402 -342 442 -341
rect 406 -346 442 -342
rect 672 -341 682 -340
rect 672 -345 678 -341
rect 260 -350 286 -346
rect 85 -356 101 -352
rect 85 -357 105 -356
rect -30 -361 -20 -360
rect -30 -365 -24 -361
rect 85 -365 105 -359
rect 256 -359 272 -355
rect 256 -360 276 -359
rect 570 -356 576 -352
rect 566 -357 576 -356
rect 672 -353 678 -349
rect 672 -354 682 -353
rect -30 -373 -24 -369
rect 85 -368 105 -367
rect 89 -372 105 -368
rect 256 -368 276 -362
rect 566 -360 576 -359
rect 566 -364 572 -360
rect 672 -362 682 -356
rect 672 -365 682 -364
rect 676 -369 682 -365
rect -30 -374 -20 -373
rect -30 -382 -20 -376
rect 256 -371 276 -370
rect 260 -375 276 -371
rect 566 -373 572 -369
rect 566 -374 576 -373
rect 566 -377 576 -376
rect 570 -381 576 -377
rect 676 -377 682 -373
rect 672 -378 682 -377
rect -30 -385 -20 -384
rect -26 -389 -20 -385
rect 94 -388 100 -384
rect 672 -381 682 -380
rect 672 -385 678 -381
rect 90 -389 100 -388
rect -26 -397 -20 -393
rect 90 -392 100 -391
rect 90 -396 96 -392
rect -30 -398 -20 -397
rect 565 -397 581 -393
rect 676 -394 682 -390
rect 672 -395 682 -394
rect 561 -398 581 -397
rect -30 -401 -20 -400
rect -30 -405 -24 -401
rect 99 -407 105 -403
rect 256 -402 312 -398
rect 256 -403 316 -402
rect 95 -408 105 -407
rect -26 -414 -20 -410
rect -30 -415 -20 -414
rect 95 -411 105 -410
rect 95 -415 101 -411
rect 256 -411 316 -405
rect 561 -406 581 -400
rect 672 -398 682 -397
rect 672 -402 678 -398
rect -30 -418 -20 -417
rect -30 -422 -24 -418
rect -26 -430 -20 -426
rect 91 -424 107 -420
rect 256 -419 316 -413
rect 561 -409 581 -408
rect 561 -413 577 -409
rect 676 -410 682 -406
rect 672 -411 682 -410
rect 561 -414 581 -413
rect 87 -425 107 -424
rect -30 -431 -20 -430
rect -30 -439 -20 -433
rect 87 -433 107 -427
rect 256 -427 316 -421
rect 561 -422 581 -416
rect 672 -419 682 -413
rect 561 -425 581 -424
rect 565 -429 581 -425
rect 672 -422 682 -421
rect 672 -426 678 -422
rect 87 -436 107 -435
rect 87 -440 103 -436
rect 256 -435 316 -429
rect -30 -442 -20 -441
rect -30 -446 -24 -442
rect 256 -443 316 -437
rect 672 -434 678 -430
rect 672 -435 682 -434
rect -30 -454 -24 -450
rect 90 -450 96 -446
rect 256 -446 316 -445
rect 260 -450 316 -446
rect 570 -445 576 -441
rect 566 -446 576 -445
rect 672 -443 682 -437
rect 672 -446 682 -445
rect 90 -451 100 -450
rect 566 -449 576 -448
rect 566 -453 572 -449
rect 676 -450 682 -446
rect -30 -455 -20 -454
rect -30 -463 -20 -457
rect 90 -454 100 -453
rect 94 -458 100 -454
rect -30 -466 -20 -465
rect 256 -459 302 -455
rect 256 -460 306 -459
rect 676 -458 682 -454
rect 672 -459 682 -458
rect -26 -470 -20 -466
rect -26 -478 -20 -474
rect 89 -474 105 -470
rect 256 -468 306 -462
rect 672 -462 682 -461
rect 672 -466 678 -462
rect 85 -475 105 -474
rect -30 -479 -20 -478
rect -30 -482 -20 -481
rect -30 -486 -24 -482
rect 85 -483 105 -477
rect 256 -476 306 -470
rect -26 -495 -20 -491
rect 85 -486 105 -485
rect 85 -490 101 -486
rect 256 -484 306 -478
rect 85 -491 105 -490
rect -30 -496 -20 -495
rect -30 -499 -20 -498
rect -30 -503 -24 -499
rect 85 -499 105 -493
rect 256 -492 306 -486
rect 256 -495 306 -494
rect 260 -499 306 -495
rect 85 -502 105 -501
rect 89 -506 105 -502
rect -26 -511 -20 -507
rect -30 -512 -20 -511
rect -30 -520 -20 -514
rect 256 -508 292 -504
rect 256 -509 296 -508
rect -30 -523 -20 -522
rect -30 -527 -24 -523
rect 94 -522 100 -518
rect 256 -517 296 -511
rect 405 -512 461 -508
rect 405 -513 465 -512
rect 90 -523 100 -522
rect 90 -526 100 -525
rect 90 -530 96 -526
rect 256 -525 296 -519
rect 405 -521 465 -515
rect -30 -535 -24 -531
rect -30 -536 -20 -535
rect -30 -544 -20 -538
rect 256 -533 296 -527
rect 405 -529 465 -523
rect 256 -536 296 -535
rect 260 -540 296 -536
rect 405 -537 465 -531
rect -30 -547 -20 -546
rect -26 -551 -20 -547
rect 256 -549 282 -545
rect 405 -545 465 -539
rect 256 -550 286 -549
rect -26 -559 -20 -555
rect -30 -560 -20 -559
rect 256 -558 286 -552
rect 405 -553 465 -547
rect 405 -556 465 -555
rect 409 -560 465 -556
rect -30 -563 -20 -562
rect -30 -567 -24 -563
rect 256 -566 286 -560
rect -26 -576 -20 -572
rect 256 -569 286 -568
rect 260 -573 286 -569
rect -30 -577 -20 -576
rect -30 -580 -20 -579
rect -30 -584 -24 -580
rect 256 -582 272 -578
rect 256 -583 276 -582
rect -26 -592 -20 -588
rect -30 -593 -20 -592
rect -30 -601 -20 -595
rect 256 -591 276 -585
rect 256 -594 276 -593
rect 260 -598 276 -594
rect -30 -604 -20 -603
rect -30 -608 -24 -604
rect -30 -616 -24 -612
rect -30 -617 -20 -616
rect -30 -625 -20 -619
rect -30 -628 -20 -627
rect -26 -632 -20 -628
rect -26 -640 -20 -636
rect -30 -641 -20 -640
rect -30 -644 -20 -643
rect -30 -648 -24 -644
<< pdiffusion >>
rect -68 151 -52 155
rect -68 150 -48 151
rect -68 147 -48 148
rect -64 143 -48 147
rect 286 145 291 161
rect 290 141 291 145
rect 293 157 294 161
rect 293 141 298 157
rect 310 145 315 161
rect 314 141 315 145
rect 317 157 318 161
rect 317 141 322 157
rect 326 145 331 161
rect 330 141 331 145
rect 333 157 334 161
rect 333 141 338 157
rect 342 145 347 161
rect 346 141 347 145
rect 349 141 355 161
rect 357 157 358 161
rect 357 141 362 157
rect -68 127 -52 131
rect -68 126 -48 127
rect 28 126 44 130
rect 28 125 48 126
rect -68 123 -48 124
rect -64 119 -48 123
rect 28 122 48 123
rect 32 118 48 122
rect -68 111 -52 115
rect -68 110 -48 111
rect -68 107 -48 108
rect -64 103 -48 107
rect 32 109 48 113
rect 28 108 48 109
rect 28 105 48 106
rect 28 101 44 105
rect -68 95 -52 99
rect 28 100 48 101
rect 28 97 48 98
rect -68 94 -48 95
rect 32 93 48 97
rect -68 86 -48 92
rect -68 83 -48 84
rect -64 79 -48 83
rect 32 83 48 87
rect 28 82 48 83
rect 28 79 48 80
rect 28 75 44 79
rect -68 70 -52 74
rect -68 69 -48 70
rect -68 66 -48 67
rect -64 62 -48 66
rect 33 59 69 63
rect 29 58 69 59
rect 29 55 69 56
rect -68 46 -52 50
rect -68 45 -48 46
rect 29 51 65 55
rect 29 50 69 51
rect -68 42 -48 43
rect -64 38 -48 42
rect 29 42 69 48
rect 29 39 69 40
rect 29 35 65 39
rect -68 30 -52 34
rect -68 29 -48 30
rect 29 34 69 35
rect 29 31 69 32
rect -68 26 -48 27
rect -64 22 -48 26
rect 33 27 69 31
rect -68 14 -52 18
rect -68 13 -48 14
rect 28 11 44 15
rect -68 5 -48 11
rect 28 10 48 11
rect 634 11 650 15
rect 634 10 654 11
rect 28 7 48 8
rect 32 3 48 7
rect 634 7 654 8
rect -68 2 -48 3
rect -64 -2 -48 2
rect 225 0 241 4
rect 28 -6 44 -2
rect -68 -10 -52 -6
rect -68 -11 -48 -10
rect 28 -7 48 -6
rect 221 -1 241 0
rect 638 3 654 7
rect 221 -4 241 -3
rect 221 -8 237 -4
rect 28 -10 48 -9
rect -68 -14 -48 -13
rect -64 -18 -48 -14
rect 32 -14 48 -10
rect 221 -9 241 -8
rect 371 -4 387 0
rect 367 -5 387 -4
rect 367 -8 387 -7
rect 221 -12 241 -11
rect 225 -16 241 -12
rect 367 -12 383 -8
rect 367 -13 387 -12
rect 634 -13 650 -9
rect 367 -16 387 -15
rect 32 -23 48 -19
rect -68 -34 -52 -30
rect -68 -35 -48 -34
rect 28 -24 48 -23
rect 371 -20 387 -16
rect 508 -17 524 -13
rect 504 -18 524 -17
rect 634 -14 654 -13
rect 634 -17 654 -16
rect 504 -21 524 -20
rect 504 -25 520 -21
rect 638 -21 654 -17
rect 28 -27 48 -26
rect 28 -31 44 -27
rect 28 -32 48 -31
rect 634 -29 650 -25
rect 28 -35 48 -34
rect -68 -38 -48 -37
rect -64 -42 -48 -38
rect 32 -39 48 -35
rect 634 -30 654 -29
rect 634 -33 654 -32
rect 638 -37 654 -33
rect 221 -43 237 -39
rect -68 -50 -52 -46
rect -68 -51 -48 -50
rect 32 -49 48 -45
rect -68 -54 -48 -53
rect -64 -58 -48 -54
rect 28 -50 48 -49
rect 221 -44 241 -43
rect 509 -41 545 -37
rect 505 -42 545 -41
rect 505 -45 545 -44
rect 221 -47 241 -46
rect 225 -51 241 -47
rect 28 -53 48 -52
rect 28 -57 44 -53
rect 221 -52 241 -51
rect 505 -49 541 -45
rect 505 -50 545 -49
rect 634 -45 650 -41
rect 634 -46 654 -45
rect 221 -55 241 -54
rect 221 -59 237 -55
rect -68 -66 -52 -62
rect 221 -60 241 -59
rect 505 -58 545 -52
rect 634 -54 654 -48
rect 634 -57 654 -56
rect 505 -61 545 -60
rect 221 -63 241 -62
rect -68 -67 -48 -66
rect 225 -67 241 -63
rect 367 -67 383 -63
rect -68 -75 -48 -69
rect 33 -73 69 -69
rect 29 -74 69 -73
rect 367 -68 387 -67
rect 505 -65 541 -61
rect 505 -66 545 -65
rect 638 -61 654 -57
rect 505 -69 545 -68
rect 367 -71 387 -70
rect 29 -77 69 -76
rect -68 -78 -48 -77
rect -64 -82 -48 -78
rect 29 -81 65 -77
rect 29 -82 69 -81
rect 225 -76 241 -72
rect 221 -77 241 -76
rect 371 -75 387 -71
rect 367 -76 387 -75
rect 509 -73 545 -69
rect 634 -70 650 -66
rect 634 -71 654 -70
rect 634 -74 654 -73
rect 638 -78 654 -74
rect 367 -79 387 -78
rect 221 -80 241 -79
rect -68 -91 -52 -87
rect -68 -92 -48 -91
rect 29 -90 69 -84
rect 221 -84 237 -80
rect 221 -85 241 -84
rect 367 -83 383 -79
rect 367 -84 387 -83
rect 367 -87 387 -86
rect 221 -88 241 -87
rect 225 -92 241 -88
rect 371 -91 387 -87
rect 504 -89 520 -85
rect 29 -93 69 -92
rect -68 -95 -48 -94
rect -64 -99 -48 -95
rect 29 -97 65 -93
rect 29 -98 69 -97
rect 504 -90 524 -89
rect 504 -93 524 -92
rect 508 -97 524 -93
rect 634 -94 650 -90
rect 634 -95 654 -94
rect 634 -98 654 -97
rect 29 -101 69 -100
rect 33 -105 69 -101
rect 638 -102 654 -98
rect 508 -107 524 -103
rect -68 -115 -52 -111
rect -68 -116 -48 -115
rect 504 -108 524 -107
rect 634 -110 650 -106
rect 504 -111 524 -110
rect 504 -115 520 -111
rect 634 -111 654 -110
rect 634 -114 654 -113
rect -68 -119 -48 -118
rect -64 -123 -48 -119
rect 28 -121 44 -117
rect 28 -122 48 -121
rect 225 -119 241 -115
rect 221 -120 241 -119
rect 638 -118 654 -114
rect 221 -123 241 -122
rect 28 -125 48 -124
rect -68 -131 -52 -127
rect -68 -132 -48 -131
rect 32 -129 48 -125
rect 221 -127 237 -123
rect 221 -128 241 -127
rect 634 -126 650 -122
rect 221 -131 241 -130
rect -68 -135 -48 -134
rect -64 -139 -48 -135
rect 225 -135 241 -131
rect 28 -141 44 -137
rect 28 -142 48 -141
rect 221 -136 241 -135
rect 509 -131 545 -127
rect 505 -132 545 -131
rect 634 -127 654 -126
rect 505 -135 545 -134
rect 221 -139 241 -138
rect -68 -147 -52 -143
rect 221 -143 237 -139
rect 28 -145 48 -144
rect -68 -148 -48 -147
rect 32 -149 48 -145
rect 221 -144 241 -143
rect 505 -139 541 -135
rect 505 -140 545 -139
rect 634 -135 654 -129
rect 634 -138 654 -137
rect 221 -147 241 -146
rect -68 -156 -48 -150
rect 225 -151 241 -147
rect 505 -148 545 -142
rect 638 -142 654 -138
rect 505 -151 545 -150
rect 32 -158 48 -154
rect -68 -159 -48 -158
rect -64 -163 -48 -159
rect 28 -159 48 -158
rect 505 -155 541 -151
rect 221 -160 237 -156
rect 28 -162 48 -161
rect 28 -166 44 -162
rect -68 -172 -52 -168
rect -68 -173 -48 -172
rect 28 -167 48 -166
rect 221 -161 241 -160
rect 505 -156 545 -155
rect 634 -151 650 -147
rect 634 -152 654 -151
rect 634 -155 654 -154
rect 505 -159 545 -158
rect 221 -164 241 -163
rect 225 -168 241 -164
rect 28 -170 48 -169
rect 32 -174 48 -170
rect 221 -169 241 -168
rect 371 -164 387 -160
rect 367 -165 387 -164
rect 509 -163 545 -159
rect 638 -159 654 -155
rect 367 -168 387 -167
rect 221 -172 241 -171
rect -68 -176 -48 -175
rect -64 -180 -48 -176
rect 221 -176 237 -172
rect 221 -177 241 -176
rect 367 -172 383 -168
rect 367 -173 387 -172
rect 634 -175 650 -171
rect 367 -176 387 -175
rect 221 -180 241 -179
rect 32 -184 48 -180
rect 28 -185 48 -184
rect 225 -184 241 -180
rect 371 -180 387 -176
rect 367 -181 387 -180
rect 504 -179 520 -175
rect 504 -180 524 -179
rect 634 -176 654 -175
rect 634 -179 654 -178
rect 504 -183 524 -182
rect 367 -184 387 -183
rect 28 -188 48 -187
rect -68 -196 -52 -192
rect -68 -197 -48 -196
rect 28 -192 44 -188
rect 367 -188 383 -184
rect -68 -200 -48 -199
rect -64 -204 -48 -200
rect 225 -193 241 -189
rect 221 -194 241 -193
rect 367 -189 387 -188
rect 508 -187 524 -183
rect 638 -183 654 -179
rect 634 -191 650 -187
rect 367 -192 387 -191
rect 371 -196 387 -192
rect 508 -196 524 -192
rect 221 -197 241 -196
rect 221 -201 237 -197
rect 33 -208 69 -204
rect -68 -212 -52 -208
rect -68 -213 -48 -212
rect 29 -209 69 -208
rect 221 -202 241 -201
rect 504 -197 524 -196
rect 634 -192 654 -191
rect 634 -195 654 -194
rect 638 -199 654 -195
rect 504 -200 524 -199
rect 504 -204 520 -200
rect 221 -205 241 -204
rect 29 -212 69 -211
rect -68 -216 -48 -215
rect -64 -220 -48 -216
rect 29 -216 65 -212
rect 29 -217 69 -216
rect 225 -209 241 -205
rect 634 -207 650 -203
rect 634 -208 654 -207
rect -68 -228 -52 -224
rect 29 -225 69 -219
rect 509 -220 545 -216
rect 505 -221 545 -220
rect 634 -216 654 -210
rect 634 -219 654 -218
rect 505 -224 545 -223
rect 29 -228 69 -227
rect -68 -229 -48 -228
rect -68 -237 -48 -231
rect 29 -232 65 -228
rect 29 -233 69 -232
rect 505 -228 541 -224
rect 505 -229 545 -228
rect 638 -223 654 -219
rect 29 -236 69 -235
rect -68 -240 -48 -239
rect -64 -244 -48 -240
rect 33 -240 69 -236
rect 221 -236 237 -232
rect 221 -237 241 -236
rect 221 -240 241 -239
rect 225 -244 241 -240
rect 221 -245 241 -244
rect 505 -237 545 -231
rect 634 -232 650 -228
rect 634 -233 654 -232
rect 634 -236 654 -235
rect 505 -240 545 -239
rect 505 -244 541 -240
rect 221 -248 241 -247
rect -68 -253 -52 -249
rect -68 -254 -48 -253
rect 221 -252 237 -248
rect 28 -256 44 -252
rect -68 -257 -48 -256
rect -64 -261 -48 -257
rect 28 -257 48 -256
rect 221 -253 241 -252
rect 505 -245 545 -244
rect 638 -240 654 -236
rect 505 -248 545 -247
rect 509 -252 545 -248
rect 221 -256 241 -255
rect 28 -260 48 -259
rect 32 -264 48 -260
rect 225 -260 241 -256
rect 221 -261 241 -260
rect 634 -256 650 -252
rect 634 -257 654 -256
rect 634 -260 654 -259
rect 221 -264 241 -263
rect 221 -268 237 -264
rect -68 -277 -52 -273
rect -68 -278 -48 -277
rect 28 -273 44 -269
rect 28 -274 48 -273
rect 221 -269 241 -268
rect 638 -264 654 -260
rect 504 -268 520 -264
rect 221 -272 241 -271
rect 225 -276 241 -272
rect 504 -269 524 -268
rect 504 -272 524 -271
rect 508 -276 524 -272
rect 634 -272 650 -268
rect 634 -273 654 -272
rect 634 -276 654 -275
rect 28 -277 48 -276
rect -68 -281 -48 -280
rect -64 -285 -48 -281
rect 32 -281 48 -277
rect 638 -280 654 -276
rect -68 -293 -52 -289
rect -68 -294 -48 -293
rect 32 -290 48 -286
rect -68 -297 -48 -296
rect -64 -301 -48 -297
rect 28 -291 48 -290
rect 225 -285 241 -281
rect 221 -286 241 -285
rect 508 -284 524 -280
rect 504 -285 524 -284
rect 504 -288 524 -287
rect 221 -289 241 -288
rect 221 -293 237 -289
rect 28 -294 48 -293
rect 28 -298 44 -294
rect 28 -299 48 -298
rect 221 -294 241 -293
rect 504 -292 520 -288
rect 634 -288 650 -284
rect 634 -289 654 -288
rect 221 -297 241 -296
rect 28 -302 48 -301
rect -68 -309 -52 -305
rect 32 -306 48 -302
rect 225 -301 241 -297
rect 221 -302 241 -301
rect 634 -297 654 -291
rect 634 -300 654 -299
rect 221 -305 241 -304
rect 221 -309 237 -305
rect -68 -310 -48 -309
rect -68 -318 -48 -312
rect 32 -316 48 -312
rect 28 -317 48 -316
rect 221 -310 241 -309
rect 368 -306 384 -302
rect 368 -307 388 -306
rect 638 -304 654 -300
rect 509 -308 545 -304
rect 505 -309 545 -308
rect 368 -310 388 -309
rect 221 -313 241 -312
rect 225 -317 241 -313
rect 372 -314 388 -310
rect 368 -315 388 -314
rect 505 -312 545 -311
rect 505 -316 541 -312
rect 505 -317 545 -316
rect 634 -313 650 -309
rect 634 -314 654 -313
rect 368 -318 388 -317
rect 28 -320 48 -319
rect -68 -321 -48 -320
rect -64 -325 -48 -321
rect 28 -324 44 -320
rect 368 -322 384 -318
rect 221 -326 237 -322
rect -68 -333 -52 -329
rect -68 -334 -48 -333
rect 221 -327 241 -326
rect 368 -323 388 -322
rect 368 -326 388 -325
rect 221 -330 241 -329
rect 225 -334 241 -330
rect -68 -337 -48 -336
rect -64 -341 -48 -337
rect 33 -340 69 -336
rect 29 -341 69 -340
rect 221 -335 241 -334
rect 372 -330 388 -326
rect 368 -331 388 -330
rect 505 -325 545 -319
rect 634 -317 654 -316
rect 638 -321 654 -317
rect 505 -328 545 -327
rect 505 -332 541 -328
rect 368 -334 388 -333
rect 221 -338 241 -337
rect 29 -344 69 -343
rect 29 -348 65 -344
rect 29 -349 69 -348
rect 221 -342 237 -338
rect 221 -343 241 -342
rect 368 -338 384 -334
rect 368 -339 388 -338
rect 505 -333 545 -332
rect 505 -336 545 -335
rect 509 -340 545 -336
rect 634 -337 650 -333
rect 634 -338 654 -337
rect 634 -341 654 -340
rect 368 -342 388 -341
rect 221 -346 241 -345
rect -68 -357 -52 -353
rect -68 -358 -48 -357
rect 29 -357 69 -351
rect 225 -350 241 -346
rect 372 -346 388 -342
rect 638 -345 654 -341
rect 225 -359 241 -355
rect 29 -360 69 -359
rect -68 -361 -48 -360
rect -64 -365 -48 -361
rect 29 -364 65 -360
rect 29 -365 69 -364
rect 221 -360 241 -359
rect 504 -356 520 -352
rect 504 -357 524 -356
rect 634 -353 650 -349
rect 634 -354 654 -353
rect 634 -357 654 -356
rect 504 -360 524 -359
rect 221 -363 241 -362
rect 221 -367 237 -363
rect 29 -368 69 -367
rect -68 -373 -52 -369
rect -68 -374 -48 -373
rect 33 -372 69 -368
rect 221 -368 241 -367
rect 508 -364 524 -360
rect 638 -361 654 -357
rect 634 -369 650 -365
rect 221 -371 241 -370
rect -68 -377 -48 -376
rect -64 -381 -48 -377
rect 225 -375 241 -371
rect 508 -373 524 -369
rect 504 -374 524 -373
rect 634 -370 654 -369
rect 504 -377 524 -376
rect 504 -381 520 -377
rect 634 -378 654 -372
rect 634 -381 654 -380
rect -68 -389 -52 -385
rect 28 -388 44 -384
rect -68 -390 -48 -389
rect 28 -389 48 -388
rect 638 -385 654 -381
rect 28 -392 48 -391
rect -68 -398 -48 -392
rect 32 -396 48 -392
rect 509 -397 545 -393
rect 505 -398 545 -397
rect 634 -394 650 -390
rect 634 -395 654 -394
rect -68 -401 -48 -400
rect -64 -405 -48 -401
rect 225 -402 241 -398
rect 28 -407 44 -403
rect 28 -408 48 -407
rect 221 -403 241 -402
rect 505 -401 545 -400
rect 505 -405 541 -401
rect 221 -406 241 -405
rect 221 -410 237 -406
rect -68 -414 -52 -410
rect -68 -415 -48 -414
rect 28 -411 48 -410
rect 32 -415 48 -411
rect 221 -411 241 -410
rect 505 -406 545 -405
rect 634 -398 654 -397
rect 638 -402 654 -398
rect 221 -414 241 -413
rect -68 -418 -48 -417
rect -64 -422 -48 -418
rect 225 -418 241 -414
rect 32 -424 48 -420
rect 28 -425 48 -424
rect 221 -419 241 -418
rect 505 -414 545 -408
rect 505 -417 545 -416
rect 505 -421 541 -417
rect 221 -422 241 -421
rect 221 -426 237 -422
rect 28 -428 48 -427
rect -68 -438 -52 -434
rect -68 -439 -48 -438
rect 28 -432 44 -428
rect 28 -433 48 -432
rect 221 -427 241 -426
rect 505 -422 545 -421
rect 634 -418 650 -414
rect 634 -419 654 -418
rect 634 -422 654 -421
rect 505 -425 545 -424
rect 509 -429 545 -425
rect 638 -426 654 -422
rect 221 -430 241 -429
rect 225 -434 241 -430
rect 28 -436 48 -435
rect 32 -440 48 -436
rect 221 -435 241 -434
rect 634 -434 650 -430
rect 221 -438 241 -437
rect -68 -442 -48 -441
rect -64 -446 -48 -442
rect 221 -442 237 -438
rect 221 -443 241 -442
rect 634 -435 654 -434
rect 634 -438 654 -437
rect 504 -445 520 -441
rect 221 -446 241 -445
rect 32 -450 48 -446
rect -68 -454 -52 -450
rect -68 -455 -48 -454
rect 28 -451 48 -450
rect 225 -450 241 -446
rect 504 -446 524 -445
rect 638 -442 654 -438
rect 504 -449 524 -448
rect 508 -453 524 -449
rect 634 -450 650 -446
rect 28 -454 48 -453
rect -68 -458 -48 -457
rect -64 -462 -48 -458
rect 28 -458 44 -454
rect 634 -451 654 -450
rect 221 -459 237 -455
rect 221 -460 241 -459
rect 634 -459 654 -453
rect 634 -462 654 -461
rect 221 -463 241 -462
rect -68 -470 -52 -466
rect 225 -467 241 -463
rect -68 -471 -48 -470
rect -68 -479 -48 -473
rect 33 -474 69 -470
rect 29 -475 69 -474
rect 221 -468 241 -467
rect 638 -466 654 -462
rect 221 -471 241 -470
rect 29 -478 69 -477
rect -68 -482 -48 -481
rect -64 -486 -48 -482
rect 29 -482 65 -478
rect 29 -483 69 -482
rect 221 -475 237 -471
rect 221 -476 241 -475
rect 221 -479 241 -478
rect -68 -495 -52 -491
rect -68 -496 -48 -495
rect 29 -491 69 -485
rect 225 -483 241 -479
rect 221 -484 241 -483
rect 221 -487 241 -486
rect 221 -491 237 -487
rect 29 -494 69 -493
rect 29 -498 65 -494
rect -68 -499 -48 -498
rect -64 -503 -48 -499
rect 29 -499 69 -498
rect 221 -492 241 -491
rect 221 -495 241 -494
rect 225 -499 241 -495
rect 29 -502 69 -501
rect 33 -506 69 -502
rect 225 -508 241 -504
rect -68 -519 -52 -515
rect -68 -520 -48 -519
rect 221 -509 241 -508
rect 221 -512 241 -511
rect 221 -516 237 -512
rect 28 -522 44 -518
rect -68 -523 -48 -522
rect -64 -527 -48 -523
rect 28 -523 48 -522
rect 221 -517 241 -516
rect 372 -512 388 -508
rect 368 -513 388 -512
rect 368 -516 388 -515
rect 221 -520 241 -519
rect 225 -524 241 -520
rect 28 -526 48 -525
rect 32 -530 48 -526
rect 221 -525 241 -524
rect 368 -520 384 -516
rect 368 -521 388 -520
rect 368 -524 388 -523
rect 221 -528 241 -527
rect -68 -535 -52 -531
rect -68 -536 -48 -535
rect 221 -532 237 -528
rect -68 -539 -48 -538
rect -64 -543 -48 -539
rect 221 -533 241 -532
rect 372 -528 388 -524
rect 368 -529 388 -528
rect 368 -532 388 -531
rect 221 -536 241 -535
rect 225 -540 241 -536
rect 368 -536 384 -532
rect 368 -537 388 -536
rect 368 -540 388 -539
rect 372 -544 388 -540
rect -68 -551 -52 -547
rect 221 -549 237 -545
rect -68 -552 -48 -551
rect 221 -550 241 -549
rect 368 -545 388 -544
rect 368 -548 388 -547
rect 368 -552 384 -548
rect 221 -553 241 -552
rect -68 -560 -48 -554
rect 225 -557 241 -553
rect 221 -558 241 -557
rect 368 -553 388 -552
rect 368 -556 388 -555
rect 372 -560 388 -556
rect 221 -561 241 -560
rect -68 -563 -48 -562
rect -64 -567 -48 -563
rect 221 -565 237 -561
rect 221 -566 241 -565
rect 221 -569 241 -568
rect -68 -576 -52 -572
rect -68 -577 -48 -576
rect 225 -573 241 -569
rect -68 -580 -48 -579
rect -64 -584 -48 -580
rect 225 -582 241 -578
rect 221 -583 241 -582
rect 221 -586 241 -585
rect 221 -590 237 -586
rect -68 -600 -52 -596
rect -68 -601 -48 -600
rect 221 -591 241 -590
rect 221 -594 241 -593
rect 225 -598 241 -594
rect -68 -604 -48 -603
rect -64 -608 -48 -604
rect -68 -616 -52 -612
rect -68 -617 -48 -616
rect -68 -620 -48 -619
rect -64 -624 -48 -620
rect -68 -632 -52 -628
rect -68 -633 -48 -632
rect -68 -641 -48 -635
rect -68 -644 -48 -643
rect -64 -648 -48 -644
<< ndcontact >>
rect -30 151 -26 155
rect -24 143 -20 147
rect -30 135 -26 139
rect 95 126 99 130
rect -24 119 -20 123
rect 101 118 105 122
rect 286 119 290 123
rect -24 111 -20 115
rect 294 113 298 117
rect 302 119 306 123
rect 318 113 322 117
rect 326 113 330 117
rect 342 119 346 123
rect 350 119 354 123
rect 358 113 362 117
rect 87 109 91 113
rect -30 95 -26 99
rect 103 93 107 97
rect -30 87 -26 91
rect -24 79 -20 83
rect 96 83 100 87
rect 90 75 94 79
rect -30 70 -26 74
rect -24 62 -20 66
rect 85 59 89 63
rect -30 54 -26 58
rect -24 38 -20 42
rect 101 43 105 47
rect -24 30 -20 34
rect 85 27 89 31
rect -30 14 -26 18
rect -30 6 -26 10
rect 90 11 94 15
rect 672 11 676 15
rect 96 3 100 7
rect -24 -2 -20 2
rect -30 -10 -26 -6
rect 95 -6 99 -2
rect 273 0 277 4
rect 678 3 682 7
rect 101 -14 105 -10
rect 417 -4 421 0
rect 672 -5 676 -1
rect -24 -18 -20 -14
rect 257 -16 261 -12
rect -30 -26 -26 -22
rect 87 -23 91 -19
rect 401 -20 405 -16
rect 572 -17 576 -13
rect 678 -21 682 -17
rect 566 -25 570 -21
rect -24 -42 -20 -38
rect 678 -29 682 -25
rect 103 -39 107 -35
rect -24 -50 -20 -46
rect 96 -49 100 -45
rect 283 -43 287 -39
rect 561 -41 565 -37
rect 90 -57 94 -53
rect 672 -45 676 -41
rect -30 -66 -26 -62
rect 577 -57 581 -53
rect 672 -53 676 -49
rect 257 -67 261 -63
rect -30 -74 -26 -70
rect 85 -73 89 -69
rect 429 -67 433 -63
rect 678 -61 682 -57
rect -24 -82 -20 -78
rect 273 -76 277 -72
rect 561 -73 565 -69
rect 672 -70 676 -66
rect 678 -78 682 -74
rect -30 -91 -26 -87
rect 101 -89 105 -85
rect 257 -92 261 -88
rect 403 -91 407 -87
rect -24 -99 -20 -95
rect 566 -89 570 -85
rect 672 -86 676 -82
rect 572 -97 576 -93
rect -30 -107 -26 -103
rect 85 -105 89 -101
rect 678 -102 682 -98
rect 572 -107 576 -103
rect 566 -115 570 -111
rect 678 -110 682 -106
rect -24 -123 -20 -119
rect 90 -121 94 -117
rect 292 -119 296 -115
rect -24 -131 -20 -127
rect 96 -129 100 -125
rect 672 -126 676 -122
rect 95 -141 99 -137
rect 561 -131 565 -127
rect -30 -147 -26 -143
rect 101 -149 105 -145
rect 672 -134 676 -130
rect 256 -151 260 -147
rect 678 -142 682 -138
rect 577 -147 581 -143
rect -30 -155 -26 -151
rect -24 -163 -20 -159
rect 87 -158 91 -154
rect -30 -172 -26 -168
rect 282 -160 286 -156
rect 672 -151 676 -147
rect 103 -174 107 -170
rect 428 -164 432 -160
rect 678 -159 682 -155
rect 561 -163 565 -159
rect 672 -167 676 -163
rect -24 -180 -20 -176
rect -30 -188 -26 -184
rect 96 -184 100 -180
rect 256 -184 260 -180
rect 566 -179 570 -175
rect 90 -192 94 -188
rect 272 -193 276 -189
rect 678 -183 682 -179
rect 572 -187 576 -183
rect 402 -196 406 -192
rect -24 -204 -20 -200
rect -24 -212 -20 -208
rect 85 -208 89 -204
rect 572 -196 576 -192
rect 678 -191 682 -187
rect 566 -204 570 -200
rect 256 -209 260 -205
rect 672 -207 676 -203
rect -30 -228 -26 -224
rect 101 -224 105 -220
rect 561 -220 565 -216
rect 672 -215 676 -211
rect -30 -236 -26 -232
rect 678 -223 682 -219
rect 85 -240 89 -236
rect 302 -236 306 -232
rect -24 -244 -20 -240
rect 577 -236 581 -232
rect 672 -232 676 -228
rect -30 -253 -26 -249
rect -24 -261 -20 -257
rect 90 -256 94 -252
rect 678 -240 682 -236
rect 672 -248 676 -244
rect 561 -252 565 -248
rect 96 -264 100 -260
rect -30 -269 -26 -265
rect 95 -273 99 -269
rect 678 -264 682 -260
rect 566 -268 570 -264
rect 256 -276 260 -272
rect 572 -276 576 -272
rect 678 -272 682 -268
rect 101 -281 105 -277
rect -24 -285 -20 -281
rect -24 -293 -20 -289
rect 87 -290 91 -286
rect 292 -285 296 -281
rect 572 -284 576 -280
rect 672 -288 676 -284
rect 566 -292 570 -288
rect -30 -309 -26 -305
rect 103 -306 107 -302
rect 672 -296 676 -292
rect -30 -317 -26 -313
rect 96 -316 100 -312
rect 438 -306 442 -302
rect 678 -304 682 -300
rect 561 -308 565 -304
rect 256 -317 260 -313
rect 672 -313 676 -309
rect -24 -325 -20 -321
rect 90 -324 94 -320
rect -30 -333 -26 -329
rect 282 -326 286 -322
rect -24 -341 -20 -337
rect 85 -340 89 -336
rect 577 -324 581 -320
rect 678 -321 682 -317
rect -30 -349 -26 -345
rect 672 -329 676 -325
rect 561 -340 565 -336
rect 402 -346 406 -342
rect 678 -345 682 -341
rect 256 -350 260 -346
rect 101 -356 105 -352
rect -24 -365 -20 -361
rect 272 -359 276 -355
rect 566 -356 570 -352
rect 678 -353 682 -349
rect -24 -373 -20 -369
rect 85 -372 89 -368
rect 572 -364 576 -360
rect 672 -369 676 -365
rect 256 -375 260 -371
rect 572 -373 576 -369
rect 566 -381 570 -377
rect 672 -377 676 -373
rect -30 -389 -26 -385
rect 90 -388 94 -384
rect 678 -385 682 -381
rect -30 -397 -26 -393
rect 96 -396 100 -392
rect 561 -397 565 -393
rect 672 -394 676 -390
rect -24 -405 -20 -401
rect 95 -407 99 -403
rect 312 -402 316 -398
rect -30 -414 -26 -410
rect 101 -415 105 -411
rect 678 -402 682 -398
rect -24 -422 -20 -418
rect -30 -430 -26 -426
rect 87 -424 91 -420
rect 577 -413 581 -409
rect 672 -410 676 -406
rect 561 -429 565 -425
rect 678 -426 682 -422
rect 103 -440 107 -436
rect -24 -446 -20 -442
rect 678 -434 682 -430
rect -24 -454 -20 -450
rect 96 -450 100 -446
rect 256 -450 260 -446
rect 566 -445 570 -441
rect 572 -453 576 -449
rect 672 -450 676 -446
rect 90 -458 94 -454
rect 302 -459 306 -455
rect 672 -458 676 -454
rect -30 -470 -26 -466
rect -30 -478 -26 -474
rect 85 -474 89 -470
rect 678 -466 682 -462
rect -24 -486 -20 -482
rect -30 -495 -26 -491
rect 101 -490 105 -486
rect -24 -503 -20 -499
rect 256 -499 260 -495
rect 85 -506 89 -502
rect -30 -511 -26 -507
rect 292 -508 296 -504
rect -24 -527 -20 -523
rect 90 -522 94 -518
rect 461 -512 465 -508
rect 96 -530 100 -526
rect -24 -535 -20 -531
rect 256 -540 260 -536
rect -30 -551 -26 -547
rect 282 -549 286 -545
rect -30 -559 -26 -555
rect 405 -560 409 -556
rect -24 -567 -20 -563
rect -30 -576 -26 -572
rect 256 -573 260 -569
rect -24 -584 -20 -580
rect 272 -582 276 -578
rect -30 -592 -26 -588
rect 256 -598 260 -594
rect -24 -608 -20 -604
rect -24 -616 -20 -612
rect -30 -632 -26 -628
rect -30 -640 -26 -636
rect -24 -648 -20 -644
<< pdcontact >>
rect -52 151 -48 155
rect -68 143 -64 147
rect 286 141 290 145
rect 294 157 298 161
rect 310 141 314 145
rect 318 157 322 161
rect 326 141 330 145
rect 334 157 338 161
rect 342 141 346 145
rect 358 157 362 161
rect -52 127 -48 131
rect 44 126 48 130
rect -68 119 -64 123
rect 28 118 32 122
rect -52 111 -48 115
rect -68 103 -64 107
rect 28 109 32 113
rect 44 101 48 105
rect -52 95 -48 99
rect 28 93 32 97
rect -68 79 -64 83
rect 28 83 32 87
rect 44 75 48 79
rect -52 70 -48 74
rect -68 62 -64 66
rect 29 59 33 63
rect -52 46 -48 50
rect 65 51 69 55
rect -68 38 -64 42
rect 65 35 69 39
rect -52 30 -48 34
rect -68 22 -64 26
rect 29 27 33 31
rect -52 14 -48 18
rect 44 11 48 15
rect 650 11 654 15
rect 28 3 32 7
rect -68 -2 -64 2
rect 221 0 225 4
rect 44 -6 48 -2
rect -52 -10 -48 -6
rect 634 3 638 7
rect 237 -8 241 -4
rect -68 -18 -64 -14
rect 28 -14 32 -10
rect 367 -4 371 0
rect 221 -16 225 -12
rect 383 -12 387 -8
rect 650 -13 654 -9
rect 28 -23 32 -19
rect -52 -34 -48 -30
rect 367 -20 371 -16
rect 504 -17 508 -13
rect 520 -25 524 -21
rect 634 -21 638 -17
rect 44 -31 48 -27
rect 650 -29 654 -25
rect -68 -42 -64 -38
rect 28 -39 32 -35
rect 634 -37 638 -33
rect 237 -43 241 -39
rect -52 -50 -48 -46
rect 28 -49 32 -45
rect -68 -58 -64 -54
rect 505 -41 509 -37
rect 221 -51 225 -47
rect 44 -57 48 -53
rect 541 -49 545 -45
rect 650 -45 654 -41
rect 237 -59 241 -55
rect -52 -66 -48 -62
rect 221 -67 225 -63
rect 383 -67 387 -63
rect 29 -73 33 -69
rect 541 -65 545 -61
rect 634 -61 638 -57
rect -68 -82 -64 -78
rect 65 -81 69 -77
rect 221 -76 225 -72
rect 367 -75 371 -71
rect 505 -73 509 -69
rect 650 -70 654 -66
rect 634 -78 638 -74
rect -52 -91 -48 -87
rect 237 -84 241 -80
rect 383 -83 387 -79
rect 221 -92 225 -88
rect 367 -91 371 -87
rect 520 -89 524 -85
rect -68 -99 -64 -95
rect 65 -97 69 -93
rect 504 -97 508 -93
rect 650 -94 654 -90
rect 29 -105 33 -101
rect 634 -102 638 -98
rect 504 -107 508 -103
rect -52 -115 -48 -111
rect 650 -110 654 -106
rect 520 -115 524 -111
rect -68 -123 -64 -119
rect 44 -121 48 -117
rect 221 -119 225 -115
rect 634 -118 638 -114
rect -52 -131 -48 -127
rect 28 -129 32 -125
rect 237 -127 241 -123
rect 650 -126 654 -122
rect -68 -139 -64 -135
rect 221 -135 225 -131
rect 44 -141 48 -137
rect 505 -131 509 -127
rect -52 -147 -48 -143
rect 237 -143 241 -139
rect 28 -149 32 -145
rect 541 -139 545 -135
rect 221 -151 225 -147
rect 634 -142 638 -138
rect 28 -158 32 -154
rect -68 -163 -64 -159
rect 541 -155 545 -151
rect 237 -160 241 -156
rect 44 -166 48 -162
rect -52 -172 -48 -168
rect 650 -151 654 -147
rect 221 -168 225 -164
rect 28 -174 32 -170
rect 367 -164 371 -160
rect 505 -163 509 -159
rect 634 -159 638 -155
rect -68 -180 -64 -176
rect 237 -176 241 -172
rect 383 -172 387 -168
rect 650 -175 654 -171
rect 28 -184 32 -180
rect 221 -184 225 -180
rect 367 -180 371 -176
rect 520 -179 524 -175
rect -52 -196 -48 -192
rect 44 -192 48 -188
rect 383 -188 387 -184
rect -68 -204 -64 -200
rect 221 -193 225 -189
rect 504 -187 508 -183
rect 634 -183 638 -179
rect 650 -191 654 -187
rect 367 -196 371 -192
rect 504 -196 508 -192
rect 237 -201 241 -197
rect 29 -208 33 -204
rect -52 -212 -48 -208
rect 634 -199 638 -195
rect 520 -204 524 -200
rect -68 -220 -64 -216
rect 65 -216 69 -212
rect 221 -209 225 -205
rect 650 -207 654 -203
rect -52 -228 -48 -224
rect 505 -220 509 -216
rect 65 -232 69 -228
rect 541 -228 545 -224
rect 634 -223 638 -219
rect -68 -244 -64 -240
rect 29 -240 33 -236
rect 237 -236 241 -232
rect 221 -244 225 -240
rect 650 -232 654 -228
rect 541 -244 545 -240
rect -52 -253 -48 -249
rect 237 -252 241 -248
rect 44 -256 48 -252
rect -68 -261 -64 -257
rect 634 -240 638 -236
rect 505 -252 509 -248
rect 28 -264 32 -260
rect 221 -260 225 -256
rect 650 -256 654 -252
rect 237 -268 241 -264
rect -52 -277 -48 -273
rect 44 -273 48 -269
rect 634 -264 638 -260
rect 520 -268 524 -264
rect 221 -276 225 -272
rect 504 -276 508 -272
rect 650 -272 654 -268
rect -68 -285 -64 -281
rect 28 -281 32 -277
rect 634 -280 638 -276
rect -52 -293 -48 -289
rect 28 -290 32 -286
rect -68 -301 -64 -297
rect 221 -285 225 -281
rect 504 -284 508 -280
rect 237 -293 241 -289
rect 44 -298 48 -294
rect 520 -292 524 -288
rect 650 -288 654 -284
rect -52 -309 -48 -305
rect 28 -306 32 -302
rect 221 -301 225 -297
rect 237 -309 241 -305
rect 28 -316 32 -312
rect 384 -306 388 -302
rect 634 -304 638 -300
rect 505 -308 509 -304
rect 221 -317 225 -313
rect 368 -314 372 -310
rect 541 -316 545 -312
rect 650 -313 654 -309
rect -68 -325 -64 -321
rect 44 -324 48 -320
rect 384 -322 388 -318
rect 237 -326 241 -322
rect -52 -333 -48 -329
rect 221 -334 225 -330
rect -68 -341 -64 -337
rect 29 -340 33 -336
rect 368 -330 372 -326
rect 634 -321 638 -317
rect 541 -332 545 -328
rect 65 -348 69 -344
rect 237 -342 241 -338
rect 384 -338 388 -334
rect 505 -340 509 -336
rect 650 -337 654 -333
rect -52 -357 -48 -353
rect 221 -350 225 -346
rect 368 -346 372 -342
rect 634 -345 638 -341
rect 221 -359 225 -355
rect -68 -365 -64 -361
rect 65 -364 69 -360
rect 520 -356 524 -352
rect 650 -353 654 -349
rect 237 -367 241 -363
rect -52 -373 -48 -369
rect 29 -372 33 -368
rect 504 -364 508 -360
rect 634 -361 638 -357
rect 650 -369 654 -365
rect -68 -381 -64 -377
rect 221 -375 225 -371
rect 504 -373 508 -369
rect 520 -381 524 -377
rect -52 -389 -48 -385
rect 44 -388 48 -384
rect 634 -385 638 -381
rect 28 -396 32 -392
rect 505 -397 509 -393
rect 650 -394 654 -390
rect -68 -405 -64 -401
rect 221 -402 225 -398
rect 44 -407 48 -403
rect 541 -405 545 -401
rect 237 -410 241 -406
rect -52 -414 -48 -410
rect 28 -415 32 -411
rect 634 -402 638 -398
rect -68 -422 -64 -418
rect 221 -418 225 -414
rect 28 -424 32 -420
rect 541 -421 545 -417
rect 237 -426 241 -422
rect -52 -438 -48 -434
rect 44 -432 48 -428
rect 650 -418 654 -414
rect 505 -429 509 -425
rect 634 -426 638 -422
rect 221 -434 225 -430
rect 28 -440 32 -436
rect 650 -434 654 -430
rect -68 -446 -64 -442
rect 237 -442 241 -438
rect 520 -445 524 -441
rect 28 -450 32 -446
rect -52 -454 -48 -450
rect 221 -450 225 -446
rect 634 -442 638 -438
rect 504 -453 508 -449
rect 650 -450 654 -446
rect -68 -462 -64 -458
rect 44 -458 48 -454
rect 237 -459 241 -455
rect -52 -470 -48 -466
rect 221 -467 225 -463
rect 29 -474 33 -470
rect 634 -466 638 -462
rect -68 -486 -64 -482
rect 65 -482 69 -478
rect 237 -475 241 -471
rect -52 -495 -48 -491
rect 221 -483 225 -479
rect 237 -491 241 -487
rect 65 -498 69 -494
rect -68 -503 -64 -499
rect 221 -499 225 -495
rect 29 -506 33 -502
rect 221 -508 225 -504
rect -52 -519 -48 -515
rect 237 -516 241 -512
rect 44 -522 48 -518
rect -68 -527 -64 -523
rect 368 -512 372 -508
rect 221 -524 225 -520
rect 28 -530 32 -526
rect 384 -520 388 -516
rect -52 -535 -48 -531
rect 237 -532 241 -528
rect -68 -543 -64 -539
rect 368 -528 372 -524
rect 221 -540 225 -536
rect 384 -536 388 -532
rect 368 -544 372 -540
rect -52 -551 -48 -547
rect 237 -549 241 -545
rect 384 -552 388 -548
rect 221 -557 225 -553
rect 368 -560 372 -556
rect -68 -567 -64 -563
rect 237 -565 241 -561
rect -52 -576 -48 -572
rect 221 -573 225 -569
rect -68 -584 -64 -580
rect 221 -582 225 -578
rect 237 -590 241 -586
rect -52 -600 -48 -596
rect 221 -598 225 -594
rect -68 -608 -64 -604
rect -52 -616 -48 -612
rect -68 -624 -64 -620
rect -52 -632 -48 -628
rect -68 -648 -64 -644
<< psubstratepcontact >>
rect 358 104 362 108
rect -15 79 -11 83
rect 111 43 115 47
rect -15 -2 -11 2
rect 330 0 334 4
rect 472 -4 476 0
rect 587 -57 591 -53
rect 472 -67 476 -63
rect 687 -61 691 -57
rect -15 -82 -11 -78
rect 111 -89 115 -85
rect 687 -143 691 -138
rect 587 -147 591 -143
rect -15 -163 -11 -159
rect 472 -164 476 -160
rect 111 -224 115 -220
rect 687 -223 691 -219
rect -15 -244 -11 -240
rect 587 -236 591 -232
rect 472 -306 476 -302
rect 687 -305 691 -300
rect -15 -325 -11 -321
rect 587 -324 591 -320
rect 111 -356 115 -352
rect 687 -385 691 -381
rect -15 -405 -11 -401
rect 587 -413 591 -409
rect 687 -466 691 -462
rect -15 -487 -11 -482
rect 111 -490 115 -486
rect 472 -512 476 -508
rect -15 -567 -11 -563
rect -15 -648 -11 -644
<< nsubstratencontact >>
rect 302 157 306 161
rect -68 135 -64 139
rect 25 67 29 71
rect -68 54 -64 58
rect 218 8 222 12
rect 364 4 368 8
rect 634 -5 638 -1
rect -68 -26 -64 -22
rect 219 -35 223 -31
rect 501 -33 505 -29
rect 25 -65 29 -61
rect 364 -59 368 -55
rect 634 -86 638 -82
rect -68 -107 -64 -103
rect 218 -111 222 -107
rect 501 -123 505 -119
rect 364 -156 368 -152
rect 634 -167 638 -163
rect -68 -188 -64 -184
rect 25 -200 29 -196
rect 501 -212 505 -208
rect 218 -228 222 -224
rect 634 -248 638 -244
rect -68 -269 -64 -265
rect 364 -298 368 -294
rect 501 -300 505 -296
rect 25 -332 29 -328
rect -68 -349 -64 -345
rect 634 -329 638 -325
rect 501 -389 505 -385
rect 218 -394 222 -390
rect -68 -430 -64 -426
rect 634 -410 638 -406
rect 25 -466 29 -462
rect 365 -504 369 -500
rect -68 -511 -64 -507
rect -68 -592 -64 -588
<< polysilicon >>
rect 291 161 293 164
rect 315 161 317 164
rect 331 161 333 176
rect 347 161 349 176
rect 355 161 357 176
rect -71 148 -68 150
rect -48 148 -30 150
rect -20 148 -17 150
rect -33 132 -30 134
rect -20 132 -8 134
rect -71 124 -68 126
rect -48 124 -30 126
rect -20 124 -17 126
rect 25 123 28 125
rect 48 123 95 125
rect 105 123 108 125
rect 291 123 293 141
rect 307 123 309 126
rect 315 123 317 141
rect 331 123 333 141
rect 347 138 349 141
rect 339 123 341 133
rect 355 123 357 141
rect -83 108 -68 110
rect -48 108 -30 110
rect -20 108 -8 110
rect 291 110 293 113
rect 12 106 28 108
rect 48 106 87 108
rect 107 106 110 108
rect -40 100 -30 102
rect -20 100 -17 102
rect 307 101 309 113
rect 315 110 317 113
rect 331 101 333 113
rect 339 110 341 113
rect 355 110 357 113
rect 12 98 28 100
rect 48 98 87 100
rect 107 98 110 100
rect -83 92 -68 94
rect -48 92 -45 94
rect -83 84 -68 86
rect -48 84 -30 86
rect -20 84 -17 86
rect 12 80 28 82
rect 48 80 90 82
rect 100 80 103 82
rect -71 67 -68 69
rect -48 67 -30 69
rect -20 67 -17 69
rect 26 56 29 58
rect 69 56 85 58
rect 105 56 118 58
rect -33 51 -30 53
rect -20 51 -8 53
rect 26 48 29 50
rect 69 48 85 50
rect 105 48 118 50
rect -71 43 -68 45
rect -48 43 -30 45
rect -20 43 -17 45
rect 12 40 29 42
rect 69 40 85 42
rect 105 40 108 42
rect 12 32 29 34
rect 69 32 85 34
rect 105 32 108 34
rect -83 27 -68 29
rect -48 27 -30 29
rect -20 27 -8 29
rect -40 19 -30 21
rect -20 19 -17 21
rect -83 11 -68 13
rect -48 11 -45 13
rect 12 8 28 10
rect 48 8 90 10
rect 100 8 103 10
rect 631 8 634 10
rect 654 8 672 10
rect 682 8 685 10
rect -83 3 -68 5
rect -48 3 -30 5
rect -20 3 -17 5
rect 206 -3 221 -1
rect 241 -3 257 -1
rect 277 -3 280 -1
rect 25 -9 28 -7
rect 48 -9 95 -7
rect 105 -9 108 -7
rect -71 -13 -68 -11
rect -48 -13 -30 -11
rect -20 -13 -17 -11
rect 352 -7 367 -5
rect 387 -7 401 -5
rect 421 -7 424 -5
rect 206 -11 221 -9
rect 241 -11 257 -9
rect 277 -11 280 -9
rect 669 -8 672 -6
rect 682 -8 694 -6
rect 352 -15 367 -13
rect 387 -15 401 -13
rect 421 -15 424 -13
rect -33 -29 -30 -27
rect -20 -29 -8 -27
rect 631 -16 634 -14
rect 654 -16 672 -14
rect 682 -16 685 -14
rect 488 -20 504 -18
rect 524 -20 566 -18
rect 576 -20 579 -18
rect 12 -26 28 -24
rect 48 -26 87 -24
rect 107 -26 110 -24
rect 12 -34 28 -32
rect 48 -34 87 -32
rect 107 -34 110 -32
rect -71 -37 -68 -35
rect -48 -37 -30 -35
rect -20 -37 -17 -35
rect 619 -32 634 -30
rect 654 -32 672 -30
rect 682 -32 694 -30
rect -83 -53 -68 -51
rect -48 -53 -30 -51
rect -20 -53 -8 -51
rect 662 -40 672 -38
rect 682 -40 685 -38
rect 502 -44 505 -42
rect 545 -44 561 -42
rect 581 -44 594 -42
rect 206 -46 221 -44
rect 241 -46 257 -44
rect 287 -46 290 -44
rect 12 -52 28 -50
rect 48 -52 90 -50
rect 100 -52 103 -50
rect 619 -48 634 -46
rect 654 -48 657 -46
rect 502 -52 505 -50
rect 545 -52 561 -50
rect 581 -52 594 -50
rect 206 -54 221 -52
rect 241 -54 257 -52
rect 287 -54 290 -52
rect -40 -61 -30 -59
rect -20 -61 -17 -59
rect 206 -62 221 -60
rect 241 -62 257 -60
rect 287 -62 290 -60
rect 619 -56 634 -54
rect 654 -56 672 -54
rect 682 -56 685 -54
rect 488 -60 505 -58
rect 545 -60 561 -58
rect 581 -60 584 -58
rect -83 -69 -68 -67
rect -48 -69 -45 -67
rect 352 -70 367 -68
rect 387 -70 403 -68
rect 433 -70 436 -68
rect 488 -68 505 -66
rect 545 -68 561 -66
rect 581 -68 584 -66
rect -83 -77 -68 -75
rect -48 -77 -30 -75
rect -20 -77 -17 -75
rect 26 -76 29 -74
rect 69 -76 85 -74
rect 105 -76 118 -74
rect 206 -79 221 -77
rect 241 -79 257 -77
rect 277 -79 280 -77
rect 631 -73 634 -71
rect 654 -73 672 -71
rect 682 -73 685 -71
rect 352 -78 367 -76
rect 387 -78 403 -76
rect 433 -78 436 -76
rect 26 -84 29 -82
rect 69 -84 85 -82
rect 105 -84 118 -82
rect -71 -94 -68 -92
rect -48 -94 -30 -92
rect -20 -94 -17 -92
rect 206 -87 221 -85
rect 241 -87 257 -85
rect 277 -87 280 -85
rect 352 -86 367 -84
rect 387 -86 403 -84
rect 433 -86 436 -84
rect 12 -92 29 -90
rect 69 -92 85 -90
rect 105 -92 108 -90
rect 669 -89 672 -87
rect 682 -89 694 -87
rect 488 -92 504 -90
rect 524 -92 566 -90
rect 576 -92 579 -90
rect 631 -97 634 -95
rect 654 -97 672 -95
rect 682 -97 685 -95
rect 12 -100 29 -98
rect 69 -100 85 -98
rect 105 -100 108 -98
rect -33 -110 -30 -108
rect -20 -110 -8 -108
rect 488 -110 504 -108
rect 524 -110 566 -108
rect 576 -110 579 -108
rect 619 -113 634 -111
rect 654 -113 672 -111
rect 682 -113 694 -111
rect -71 -118 -68 -116
rect -48 -118 -30 -116
rect -20 -118 -17 -116
rect 12 -124 28 -122
rect 48 -124 90 -122
rect 100 -124 103 -122
rect 206 -122 221 -120
rect 241 -122 256 -120
rect 296 -122 299 -120
rect 662 -121 672 -119
rect 682 -121 685 -119
rect 206 -130 221 -128
rect 241 -130 256 -128
rect 296 -130 299 -128
rect -83 -134 -68 -132
rect -48 -134 -30 -132
rect -20 -134 -8 -132
rect -40 -142 -30 -140
rect -20 -142 -17 -140
rect 619 -129 634 -127
rect 654 -129 657 -127
rect 502 -134 505 -132
rect 545 -134 561 -132
rect 581 -134 594 -132
rect 206 -138 221 -136
rect 241 -138 256 -136
rect 296 -138 299 -136
rect 25 -144 28 -142
rect 48 -144 95 -142
rect 105 -144 108 -142
rect -83 -150 -68 -148
rect -48 -150 -45 -148
rect 619 -137 634 -135
rect 654 -137 672 -135
rect 682 -137 685 -135
rect 502 -142 505 -140
rect 545 -142 561 -140
rect 581 -142 594 -140
rect 206 -146 221 -144
rect 241 -146 256 -144
rect 296 -146 299 -144
rect 488 -150 505 -148
rect 545 -150 561 -148
rect 581 -150 584 -148
rect -83 -158 -68 -156
rect -48 -158 -30 -156
rect -20 -158 -17 -156
rect 12 -161 28 -159
rect 48 -161 87 -159
rect 107 -161 110 -159
rect 631 -154 634 -152
rect 654 -154 672 -152
rect 682 -154 685 -152
rect 488 -158 505 -156
rect 545 -158 561 -156
rect 581 -158 584 -156
rect 206 -163 221 -161
rect 241 -163 256 -161
rect 286 -163 289 -161
rect 12 -169 28 -167
rect 48 -169 87 -167
rect 107 -169 110 -167
rect -71 -175 -68 -173
rect -48 -175 -30 -173
rect -20 -175 -17 -173
rect 351 -167 367 -165
rect 387 -167 402 -165
rect 432 -167 435 -165
rect 206 -171 221 -169
rect 241 -171 256 -169
rect 286 -171 289 -169
rect 669 -170 672 -168
rect 682 -170 694 -168
rect 351 -175 367 -173
rect 387 -175 402 -173
rect 432 -175 435 -173
rect 206 -179 221 -177
rect 241 -179 256 -177
rect 286 -179 289 -177
rect 351 -183 367 -181
rect 387 -183 402 -181
rect 432 -183 435 -181
rect 631 -178 634 -176
rect 654 -178 672 -176
rect 682 -178 685 -176
rect 488 -182 504 -180
rect 524 -182 566 -180
rect 576 -182 579 -180
rect 12 -187 28 -185
rect 48 -187 90 -185
rect 100 -187 103 -185
rect -33 -191 -30 -189
rect -20 -191 -8 -189
rect -71 -199 -68 -197
rect -48 -199 -30 -197
rect -20 -199 -17 -197
rect 351 -191 367 -189
rect 387 -191 402 -189
rect 432 -191 435 -189
rect 206 -196 221 -194
rect 241 -196 256 -194
rect 276 -196 279 -194
rect 619 -194 634 -192
rect 654 -194 672 -192
rect 682 -194 694 -192
rect 488 -199 504 -197
rect 524 -199 566 -197
rect 576 -199 579 -197
rect 206 -204 221 -202
rect 241 -204 256 -202
rect 276 -204 279 -202
rect 662 -202 672 -200
rect 682 -202 685 -200
rect 26 -211 29 -209
rect 69 -211 85 -209
rect 105 -211 118 -209
rect -83 -215 -68 -213
rect -48 -215 -30 -213
rect -20 -215 -8 -213
rect 619 -210 634 -208
rect 654 -210 657 -208
rect 26 -219 29 -217
rect 69 -219 85 -217
rect 105 -219 118 -217
rect -40 -223 -30 -221
rect -20 -223 -17 -221
rect 619 -218 634 -216
rect 654 -218 672 -216
rect 682 -218 685 -216
rect 502 -223 505 -221
rect 545 -223 561 -221
rect 581 -223 594 -221
rect 12 -227 29 -225
rect 69 -227 85 -225
rect 105 -227 108 -225
rect -83 -231 -68 -229
rect -48 -231 -45 -229
rect 502 -231 505 -229
rect 545 -231 561 -229
rect 581 -231 594 -229
rect 12 -235 29 -233
rect 69 -235 85 -233
rect 105 -235 108 -233
rect -83 -239 -68 -237
rect -48 -239 -30 -237
rect -20 -239 -17 -237
rect 206 -239 221 -237
rect 241 -239 256 -237
rect 306 -239 309 -237
rect 631 -235 634 -233
rect 654 -235 672 -233
rect 682 -235 685 -233
rect 488 -239 505 -237
rect 545 -239 561 -237
rect 581 -239 584 -237
rect 206 -247 221 -245
rect 241 -247 256 -245
rect 306 -247 309 -245
rect -71 -256 -68 -254
rect -48 -256 -30 -254
rect -20 -256 -17 -254
rect 488 -247 505 -245
rect 545 -247 561 -245
rect 581 -247 584 -245
rect 669 -251 672 -249
rect 682 -251 694 -249
rect 206 -255 221 -253
rect 241 -255 256 -253
rect 306 -255 309 -253
rect 12 -259 28 -257
rect 48 -259 90 -257
rect 100 -259 103 -257
rect 631 -259 634 -257
rect 654 -259 672 -257
rect 682 -259 685 -257
rect 206 -263 221 -261
rect 241 -263 256 -261
rect 306 -263 309 -261
rect -33 -272 -30 -270
rect -20 -272 -8 -270
rect 206 -271 221 -269
rect 241 -271 256 -269
rect 306 -271 309 -269
rect 25 -276 28 -274
rect 48 -276 95 -274
rect 105 -276 108 -274
rect 488 -271 504 -269
rect 524 -271 566 -269
rect 576 -271 579 -269
rect 619 -275 634 -273
rect 654 -275 672 -273
rect 682 -275 694 -273
rect -71 -280 -68 -278
rect -48 -280 -30 -278
rect -20 -280 -17 -278
rect -83 -296 -68 -294
rect -48 -296 -30 -294
rect -20 -296 -8 -294
rect 206 -288 221 -286
rect 241 -288 256 -286
rect 296 -288 299 -286
rect 662 -283 672 -281
rect 682 -283 685 -281
rect 488 -287 504 -285
rect 524 -287 566 -285
rect 576 -287 579 -285
rect 12 -293 28 -291
rect 48 -293 87 -291
rect 107 -293 110 -291
rect 619 -291 634 -289
rect 654 -291 657 -289
rect 206 -296 221 -294
rect 241 -296 256 -294
rect 296 -296 299 -294
rect 12 -301 28 -299
rect 48 -301 87 -299
rect 107 -301 110 -299
rect -40 -304 -30 -302
rect -20 -304 -17 -302
rect 619 -299 634 -297
rect 654 -299 672 -297
rect 682 -299 685 -297
rect 206 -304 221 -302
rect 241 -304 256 -302
rect 296 -304 299 -302
rect -83 -312 -68 -310
rect -48 -312 -45 -310
rect -83 -320 -68 -318
rect -48 -320 -30 -318
rect -20 -320 -17 -318
rect 351 -309 368 -307
rect 388 -309 402 -307
rect 442 -309 445 -307
rect 206 -312 221 -310
rect 241 -312 256 -310
rect 296 -312 299 -310
rect 12 -319 28 -317
rect 48 -319 90 -317
rect 100 -319 103 -317
rect 502 -311 505 -309
rect 545 -311 561 -309
rect 581 -311 594 -309
rect 351 -317 368 -315
rect 388 -317 402 -315
rect 442 -317 445 -315
rect 631 -316 634 -314
rect 654 -316 672 -314
rect 682 -316 685 -314
rect 502 -319 505 -317
rect 545 -319 561 -317
rect 581 -319 594 -317
rect 351 -325 368 -323
rect 388 -325 402 -323
rect 442 -325 445 -323
rect 206 -329 221 -327
rect 241 -329 256 -327
rect 286 -329 289 -327
rect -71 -336 -68 -334
rect -48 -336 -30 -334
rect -20 -336 -17 -334
rect 488 -327 505 -325
rect 545 -327 561 -325
rect 581 -327 584 -325
rect 351 -333 368 -331
rect 388 -333 402 -331
rect 442 -333 445 -331
rect 206 -337 221 -335
rect 241 -337 256 -335
rect 286 -337 289 -335
rect 26 -343 29 -341
rect 69 -343 85 -341
rect 105 -343 118 -341
rect 669 -332 672 -330
rect 682 -332 694 -330
rect 488 -335 505 -333
rect 545 -335 561 -333
rect 581 -335 584 -333
rect 351 -341 368 -339
rect 388 -341 402 -339
rect 442 -341 445 -339
rect 631 -340 634 -338
rect 654 -340 672 -338
rect 682 -340 685 -338
rect 206 -345 221 -343
rect 241 -345 256 -343
rect 286 -345 289 -343
rect -33 -352 -30 -350
rect -20 -352 -8 -350
rect 26 -351 29 -349
rect 69 -351 85 -349
rect 105 -351 118 -349
rect -71 -360 -68 -358
rect -48 -360 -30 -358
rect -20 -360 -17 -358
rect 12 -359 29 -357
rect 69 -359 85 -357
rect 105 -359 108 -357
rect 619 -356 634 -354
rect 654 -356 672 -354
rect 682 -356 694 -354
rect 488 -359 504 -357
rect 524 -359 566 -357
rect 576 -359 579 -357
rect 206 -362 221 -360
rect 241 -362 256 -360
rect 276 -362 279 -360
rect 12 -367 29 -365
rect 69 -367 85 -365
rect 105 -367 108 -365
rect 662 -364 672 -362
rect 682 -364 685 -362
rect 206 -370 221 -368
rect 241 -370 256 -368
rect 276 -370 279 -368
rect -83 -376 -68 -374
rect -48 -376 -30 -374
rect -20 -376 -8 -374
rect 619 -372 634 -370
rect 654 -372 657 -370
rect 488 -376 504 -374
rect 524 -376 566 -374
rect 576 -376 579 -374
rect 619 -380 634 -378
rect 654 -380 672 -378
rect 682 -380 685 -378
rect -40 -384 -30 -382
rect -20 -384 -17 -382
rect -83 -392 -68 -390
rect -48 -392 -45 -390
rect 12 -391 28 -389
rect 48 -391 90 -389
rect 100 -391 103 -389
rect 631 -397 634 -395
rect 654 -397 672 -395
rect 682 -397 685 -395
rect -83 -400 -68 -398
rect -48 -400 -30 -398
rect -20 -400 -17 -398
rect 502 -400 505 -398
rect 545 -400 561 -398
rect 581 -400 594 -398
rect 206 -405 221 -403
rect 241 -405 256 -403
rect 316 -405 319 -403
rect 25 -410 28 -408
rect 48 -410 95 -408
rect 105 -410 108 -408
rect 502 -408 505 -406
rect 545 -408 561 -406
rect 581 -408 594 -406
rect 206 -413 221 -411
rect 241 -413 256 -411
rect 316 -413 319 -411
rect -71 -417 -68 -415
rect -48 -417 -30 -415
rect -20 -417 -17 -415
rect 669 -413 672 -411
rect 682 -413 694 -411
rect 488 -416 505 -414
rect 545 -416 561 -414
rect 581 -416 584 -414
rect 206 -421 221 -419
rect 241 -421 256 -419
rect 316 -421 319 -419
rect 12 -427 28 -425
rect 48 -427 87 -425
rect 107 -427 110 -425
rect -33 -433 -30 -431
rect -20 -433 -8 -431
rect 631 -421 634 -419
rect 654 -421 672 -419
rect 682 -421 685 -419
rect 488 -424 505 -422
rect 545 -424 561 -422
rect 581 -424 584 -422
rect 206 -429 221 -427
rect 241 -429 256 -427
rect 316 -429 319 -427
rect 12 -435 28 -433
rect 48 -435 87 -433
rect 107 -435 110 -433
rect -71 -441 -68 -439
rect -48 -441 -30 -439
rect -20 -441 -17 -439
rect 206 -437 221 -435
rect 241 -437 256 -435
rect 316 -437 319 -435
rect 619 -437 634 -435
rect 654 -437 672 -435
rect 682 -437 694 -435
rect 206 -445 221 -443
rect 241 -445 256 -443
rect 316 -445 319 -443
rect 662 -445 672 -443
rect 682 -445 685 -443
rect 488 -448 504 -446
rect 524 -448 566 -446
rect 576 -448 579 -446
rect 12 -453 28 -451
rect 48 -453 90 -451
rect 100 -453 103 -451
rect -83 -457 -68 -455
rect -48 -457 -30 -455
rect -20 -457 -8 -455
rect 619 -453 634 -451
rect 654 -453 657 -451
rect -40 -465 -30 -463
rect -20 -465 -17 -463
rect 206 -462 221 -460
rect 241 -462 256 -460
rect 306 -462 309 -460
rect 619 -461 634 -459
rect 654 -461 672 -459
rect 682 -461 685 -459
rect -83 -473 -68 -471
rect -48 -473 -45 -471
rect 206 -470 221 -468
rect 241 -470 256 -468
rect 306 -470 309 -468
rect 26 -477 29 -475
rect 69 -477 85 -475
rect 105 -477 118 -475
rect -83 -481 -68 -479
rect -48 -481 -30 -479
rect -20 -481 -17 -479
rect 206 -478 221 -476
rect 241 -478 256 -476
rect 306 -478 309 -476
rect 26 -485 29 -483
rect 69 -485 85 -483
rect 105 -485 118 -483
rect 206 -486 221 -484
rect 241 -486 256 -484
rect 306 -486 309 -484
rect 12 -493 29 -491
rect 69 -493 85 -491
rect 105 -493 108 -491
rect -71 -498 -68 -496
rect -48 -498 -30 -496
rect -20 -498 -17 -496
rect 206 -494 221 -492
rect 241 -494 256 -492
rect 306 -494 309 -492
rect 12 -501 29 -499
rect 69 -501 85 -499
rect 105 -501 108 -499
rect -33 -514 -30 -512
rect -20 -514 -8 -512
rect 206 -511 221 -509
rect 241 -511 256 -509
rect 296 -511 299 -509
rect -71 -522 -68 -520
rect -48 -522 -30 -520
rect -20 -522 -17 -520
rect 351 -515 368 -513
rect 388 -515 405 -513
rect 465 -515 468 -513
rect 206 -519 221 -517
rect 241 -519 256 -517
rect 296 -519 299 -517
rect 12 -525 28 -523
rect 48 -525 90 -523
rect 100 -525 103 -523
rect 351 -523 368 -521
rect 388 -523 405 -521
rect 465 -523 468 -521
rect 206 -527 221 -525
rect 241 -527 256 -525
rect 296 -527 299 -525
rect -83 -538 -68 -536
rect -48 -538 -30 -536
rect -20 -538 -8 -536
rect 351 -531 368 -529
rect 388 -531 405 -529
rect 465 -531 468 -529
rect 206 -535 221 -533
rect 241 -535 256 -533
rect 296 -535 299 -533
rect 351 -539 368 -537
rect 388 -539 405 -537
rect 465 -539 468 -537
rect -40 -546 -30 -544
rect -20 -546 -17 -544
rect -83 -554 -68 -552
rect -48 -554 -45 -552
rect 351 -547 368 -545
rect 388 -547 405 -545
rect 465 -547 468 -545
rect 206 -552 221 -550
rect 241 -552 256 -550
rect 286 -552 289 -550
rect -83 -562 -68 -560
rect -48 -562 -30 -560
rect -20 -562 -17 -560
rect 351 -555 368 -553
rect 388 -555 405 -553
rect 465 -555 468 -553
rect 206 -560 221 -558
rect 241 -560 256 -558
rect 286 -560 289 -558
rect 206 -568 221 -566
rect 241 -568 256 -566
rect 286 -568 289 -566
rect -71 -579 -68 -577
rect -48 -579 -30 -577
rect -20 -579 -17 -577
rect 206 -585 221 -583
rect 241 -585 256 -583
rect 276 -585 279 -583
rect -33 -595 -30 -593
rect -20 -595 -8 -593
rect 206 -593 221 -591
rect 241 -593 256 -591
rect 276 -593 279 -591
rect -71 -603 -68 -601
rect -48 -603 -30 -601
rect -20 -603 -17 -601
rect -83 -619 -68 -617
rect -48 -619 -30 -617
rect -20 -619 -8 -617
rect -40 -627 -30 -625
rect -20 -627 -17 -625
rect -83 -635 -68 -633
rect -48 -635 -45 -633
rect -83 -643 -68 -641
rect -48 -643 -30 -641
rect -20 -643 -17 -641
<< polycontact >>
rect 330 176 334 180
rect 346 176 350 180
rect 354 176 358 180
rect -39 144 -35 148
rect -8 131 -4 135
rect -38 120 -34 124
rect 293 128 297 132
rect 317 127 321 131
rect 338 133 342 137
rect 60 119 64 123
rect -87 107 -83 111
rect -44 99 -40 103
rect -8 107 -4 111
rect 8 105 12 109
rect 8 97 12 101
rect -87 91 -83 95
rect 306 97 310 101
rect 330 97 334 101
rect -87 83 -83 87
rect 8 79 12 83
rect -39 63 -35 67
rect -8 50 -4 54
rect 118 55 122 59
rect -38 39 -34 43
rect 8 39 12 43
rect 118 47 122 51
rect -87 26 -83 30
rect 8 31 12 35
rect -44 18 -40 22
rect -8 26 -4 30
rect -87 10 -83 14
rect -87 2 -83 6
rect 8 7 12 11
rect 202 -4 206 0
rect 663 4 667 8
rect -39 -17 -35 -13
rect 60 -13 64 -9
rect 202 -12 206 -8
rect 348 -8 352 -4
rect 348 -16 352 -12
rect -8 -30 -4 -26
rect 8 -27 12 -23
rect 484 -21 488 -17
rect 694 -9 698 -5
rect 664 -20 668 -16
rect 8 -35 12 -31
rect -38 -41 -34 -37
rect 615 -33 619 -29
rect -87 -54 -83 -50
rect -44 -62 -40 -58
rect -8 -54 -4 -50
rect 8 -53 12 -49
rect 202 -47 206 -43
rect 658 -41 662 -37
rect 694 -33 698 -29
rect 202 -55 206 -51
rect 594 -45 598 -41
rect 615 -49 619 -45
rect 202 -63 206 -59
rect 484 -61 488 -57
rect 594 -53 598 -49
rect 615 -57 619 -53
rect -87 -70 -83 -66
rect -87 -78 -83 -74
rect 348 -71 352 -67
rect 484 -69 488 -65
rect 118 -77 122 -73
rect 202 -80 206 -76
rect 348 -79 352 -75
rect 663 -77 667 -73
rect 8 -93 12 -89
rect 118 -85 122 -81
rect 202 -88 206 -84
rect 348 -87 352 -83
rect -39 -98 -35 -94
rect 8 -101 12 -97
rect 484 -93 488 -89
rect 694 -90 698 -86
rect 664 -101 668 -97
rect -8 -111 -4 -107
rect 484 -111 488 -107
rect 615 -114 619 -110
rect -38 -122 -34 -118
rect 8 -125 12 -121
rect 202 -123 206 -119
rect -87 -135 -83 -131
rect 202 -131 206 -127
rect 658 -122 662 -118
rect 694 -114 698 -110
rect -44 -143 -40 -139
rect -8 -135 -4 -131
rect 202 -139 206 -135
rect 615 -130 619 -126
rect -87 -151 -83 -147
rect 60 -148 64 -144
rect 202 -147 206 -143
rect 594 -135 598 -131
rect 615 -138 619 -134
rect -87 -159 -83 -155
rect 484 -151 488 -147
rect 594 -143 598 -139
rect 8 -162 12 -158
rect 8 -170 12 -166
rect 202 -164 206 -160
rect 484 -159 488 -155
rect 202 -172 206 -168
rect 347 -168 351 -164
rect 663 -158 667 -154
rect -39 -179 -35 -175
rect 202 -180 206 -176
rect 347 -176 351 -172
rect 8 -188 12 -184
rect 347 -184 351 -180
rect 484 -183 488 -179
rect 694 -171 698 -167
rect -8 -192 -4 -188
rect -38 -203 -34 -199
rect 202 -197 206 -193
rect 347 -192 351 -188
rect 664 -182 668 -178
rect -87 -216 -83 -212
rect 202 -205 206 -201
rect 484 -200 488 -196
rect 615 -195 619 -191
rect 658 -203 662 -199
rect 694 -195 698 -191
rect -44 -224 -40 -220
rect -8 -216 -4 -212
rect 118 -212 122 -208
rect 615 -211 619 -207
rect 8 -228 12 -224
rect 118 -220 122 -216
rect 615 -219 619 -215
rect -87 -232 -83 -228
rect -87 -240 -83 -236
rect 8 -236 12 -232
rect 594 -224 598 -220
rect 202 -239 206 -235
rect 202 -248 206 -244
rect 484 -240 488 -236
rect 594 -232 598 -228
rect -39 -260 -35 -256
rect 8 -260 12 -256
rect 202 -256 206 -252
rect 484 -248 488 -244
rect 663 -239 667 -235
rect 202 -264 206 -260
rect 694 -252 698 -248
rect -8 -273 -4 -269
rect 202 -272 206 -268
rect 664 -263 668 -259
rect 484 -272 488 -268
rect 615 -276 619 -272
rect -38 -284 -34 -280
rect 60 -280 64 -276
rect -87 -297 -83 -293
rect -44 -305 -40 -301
rect -8 -297 -4 -293
rect 8 -294 12 -290
rect 202 -288 206 -284
rect 484 -288 488 -284
rect 658 -284 662 -280
rect 694 -276 698 -272
rect 8 -302 12 -298
rect 202 -297 206 -293
rect 615 -292 619 -288
rect 202 -305 206 -301
rect 615 -300 619 -296
rect -87 -313 -83 -309
rect -87 -321 -83 -317
rect 8 -320 12 -316
rect 202 -313 206 -309
rect 347 -310 351 -306
rect 347 -318 351 -314
rect 594 -312 598 -308
rect 202 -330 206 -326
rect 347 -326 351 -322
rect -39 -340 -35 -336
rect 202 -338 206 -334
rect 347 -334 351 -330
rect 484 -328 488 -324
rect 594 -320 598 -316
rect 663 -320 667 -316
rect 118 -344 122 -340
rect 202 -346 206 -342
rect 347 -342 351 -338
rect 484 -336 488 -332
rect 694 -333 698 -329
rect -8 -353 -4 -349
rect 8 -360 12 -356
rect 118 -352 122 -348
rect 664 -344 668 -340
rect -38 -364 -34 -360
rect 8 -368 12 -364
rect 202 -363 206 -359
rect 484 -360 488 -356
rect 615 -357 619 -353
rect -87 -377 -83 -373
rect 202 -371 206 -367
rect 658 -365 662 -361
rect 694 -357 698 -353
rect -44 -385 -40 -381
rect -8 -377 -4 -373
rect 484 -377 488 -373
rect 615 -373 619 -369
rect 615 -381 619 -377
rect -87 -393 -83 -389
rect 8 -392 12 -388
rect -87 -401 -83 -397
rect 202 -406 206 -402
rect 60 -414 64 -410
rect 202 -414 206 -410
rect 594 -401 598 -397
rect 663 -401 667 -397
rect -39 -421 -35 -417
rect 8 -428 12 -424
rect 202 -422 206 -418
rect 484 -417 488 -413
rect 594 -409 598 -405
rect -8 -434 -4 -430
rect 8 -436 12 -432
rect 202 -430 206 -426
rect 484 -425 488 -421
rect 694 -414 698 -410
rect 664 -425 668 -421
rect 202 -438 206 -434
rect -38 -445 -34 -441
rect 202 -446 206 -442
rect 615 -438 619 -434
rect -87 -458 -83 -454
rect 8 -454 12 -450
rect 484 -449 488 -445
rect 658 -446 662 -442
rect 694 -438 698 -434
rect -44 -466 -40 -462
rect -8 -458 -4 -454
rect 615 -454 619 -450
rect 202 -463 206 -459
rect 615 -462 619 -458
rect -87 -474 -83 -470
rect -87 -482 -83 -478
rect 202 -471 206 -467
rect 118 -478 122 -474
rect 202 -479 206 -475
rect 8 -494 12 -490
rect 118 -486 122 -482
rect 202 -487 206 -483
rect -39 -502 -35 -498
rect 8 -502 12 -498
rect 202 -495 206 -491
rect -8 -515 -4 -511
rect 202 -512 206 -508
rect -38 -526 -34 -522
rect 8 -526 12 -522
rect 202 -520 206 -516
rect 347 -516 351 -512
rect 202 -528 206 -524
rect 347 -524 351 -520
rect -87 -539 -83 -535
rect -44 -547 -40 -543
rect -8 -539 -4 -535
rect 202 -536 206 -532
rect 347 -532 351 -528
rect 347 -540 351 -536
rect -87 -555 -83 -551
rect 202 -553 206 -549
rect 347 -548 351 -544
rect -87 -563 -83 -559
rect 202 -561 206 -557
rect 347 -556 351 -552
rect 202 -569 206 -565
rect -39 -583 -35 -579
rect 202 -586 206 -582
rect -8 -596 -4 -592
rect 202 -594 206 -590
rect -38 -607 -34 -603
rect -87 -620 -83 -616
rect -44 -628 -40 -624
rect -8 -620 -4 -616
rect -87 -636 -83 -632
rect -87 -644 -83 -640
<< metal1 >>
rect -97 183 -93 188
rect -97 179 286 183
rect -97 95 -93 179
rect -80 172 19 176
rect 282 173 286 179
rect 334 176 346 180
rect -80 147 -76 172
rect -37 164 12 168
rect -37 155 -33 164
rect -48 151 -30 155
rect -80 143 -68 147
rect -15 147 -11 161
rect -80 139 -76 143
rect -39 139 -35 144
rect -20 143 -11 147
rect -80 135 -68 139
rect -44 136 -30 139
rect -80 123 -76 135
rect -44 131 -41 136
rect -48 127 -41 131
rect -80 119 -68 123
rect -15 123 -11 143
rect -87 95 -83 107
rect -97 91 -87 95
rect -80 107 -76 119
rect -38 115 -34 120
rect -20 119 -11 123
rect -15 115 -11 119
rect -48 111 -34 115
rect -20 111 -11 115
rect -80 103 -68 107
rect -97 14 -93 91
rect -80 83 -76 103
rect -48 95 -40 99
rect -37 99 -34 111
rect -37 95 -30 99
rect -43 91 -40 95
rect -43 87 -30 91
rect -15 83 -11 111
rect -8 111 -4 131
rect 8 109 12 164
rect -80 79 -68 83
rect -20 79 -15 83
rect -80 66 -76 79
rect -48 70 -30 74
rect -80 62 -68 66
rect -15 66 -11 79
rect -80 58 -76 62
rect -39 58 -35 63
rect -20 62 -11 66
rect -80 54 -68 58
rect -44 55 -30 58
rect -80 42 -76 54
rect -44 50 -41 55
rect -48 46 -41 50
rect -80 38 -68 42
rect -15 42 -11 62
rect 0 105 8 109
rect 15 150 19 172
rect 280 169 376 173
rect 294 161 298 165
rect 302 161 306 165
rect 318 161 322 165
rect 334 161 338 165
rect 358 161 362 165
rect 15 146 213 150
rect 15 122 19 146
rect 48 126 95 130
rect 15 118 28 122
rect 111 122 115 137
rect 15 113 19 118
rect 60 113 64 119
rect 105 118 115 122
rect 15 109 28 113
rect 60 109 87 113
rect -87 14 -83 26
rect -97 10 -87 14
rect -80 26 -76 38
rect -38 34 -34 39
rect -20 38 -11 42
rect -15 34 -11 38
rect -48 30 -34 34
rect -20 30 -11 34
rect -80 22 -68 26
rect -97 -66 -93 10
rect -80 2 -76 22
rect -48 14 -40 18
rect -37 18 -34 30
rect -37 14 -30 18
rect -43 10 -40 14
rect -43 6 -30 10
rect -15 2 -11 30
rect -8 30 -4 50
rect 0 35 4 105
rect 8 83 12 97
rect 8 43 12 74
rect 15 97 19 109
rect 73 105 77 109
rect 48 101 77 105
rect 111 97 115 118
rect 15 93 28 97
rect 107 93 115 97
rect 15 87 19 93
rect 111 87 115 93
rect 15 83 28 87
rect 100 83 115 87
rect 15 71 19 83
rect 48 75 90 79
rect 15 67 25 71
rect 0 31 8 35
rect 8 11 12 31
rect 15 23 19 67
rect 22 59 29 63
rect 82 61 85 63
rect 78 59 85 61
rect 22 31 25 59
rect 78 55 82 59
rect 69 51 82 55
rect 69 35 75 39
rect 22 27 29 31
rect 71 23 75 35
rect 78 31 82 51
rect 111 47 115 83
rect 105 43 111 47
rect 78 27 85 31
rect 15 19 75 23
rect 15 7 19 19
rect 48 11 90 15
rect 111 7 115 43
rect -80 -2 -68 2
rect -20 -2 -15 2
rect 15 3 28 7
rect 100 3 115 7
rect 0 0 1 1
rect -80 -14 -76 -2
rect -48 -7 -39 -6
rect -34 -7 -30 -6
rect -48 -10 -30 -7
rect -80 -18 -68 -14
rect -15 -14 -11 -2
rect -80 -22 -76 -18
rect -39 -22 -35 -17
rect -20 -18 -11 -14
rect -80 -26 -68 -22
rect -44 -25 -30 -22
rect -80 -38 -76 -26
rect -44 -30 -41 -25
rect -48 -34 -41 -30
rect -80 -42 -68 -38
rect -15 -38 -11 -18
rect 0 -23 4 -6
rect 15 -10 19 3
rect 48 -6 95 -2
rect 15 -14 28 -10
rect 111 -10 115 3
rect 15 -19 19 -14
rect 60 -19 64 -13
rect 105 -14 115 -10
rect 15 -23 28 -19
rect 60 -23 87 -19
rect -87 -66 -83 -54
rect -97 -70 -87 -66
rect -80 -54 -76 -42
rect -38 -46 -34 -41
rect -20 -42 -11 -38
rect -15 -46 -11 -42
rect -48 -50 -34 -46
rect -20 -50 -11 -46
rect -80 -58 -68 -54
rect -97 -147 -93 -70
rect -80 -78 -76 -58
rect -48 -66 -40 -62
rect -37 -62 -34 -50
rect -37 -66 -30 -62
rect -43 -70 -40 -66
rect -43 -74 -30 -70
rect -15 -78 -11 -50
rect -8 -50 -4 -30
rect 0 -27 8 -23
rect -80 -82 -68 -78
rect -20 -82 -15 -78
rect -80 -95 -76 -82
rect -48 -91 -30 -87
rect -80 -99 -68 -95
rect -15 -95 -11 -82
rect -80 -103 -76 -99
rect -39 -103 -35 -98
rect -20 -99 -11 -95
rect -80 -107 -68 -103
rect -44 -106 -30 -103
rect -80 -119 -76 -107
rect -44 -111 -41 -106
rect -48 -115 -41 -111
rect -80 -123 -68 -119
rect -15 -119 -11 -99
rect 0 -97 4 -27
rect 8 -49 12 -35
rect 8 -82 12 -53
rect 8 -89 12 -87
rect 15 -35 19 -23
rect 73 -27 77 -23
rect 48 -31 77 -27
rect 111 -35 115 -14
rect 15 -39 28 -35
rect 107 -39 115 -35
rect 15 -45 19 -39
rect 111 -45 115 -39
rect 15 -49 28 -45
rect 100 -49 115 -45
rect 15 -61 19 -49
rect 48 -57 90 -53
rect 15 -65 25 -61
rect 0 -101 8 -97
rect -87 -147 -83 -135
rect -97 -151 -87 -147
rect -80 -135 -76 -123
rect -38 -127 -34 -122
rect -20 -123 -11 -119
rect -15 -127 -11 -123
rect -48 -131 -34 -127
rect -20 -131 -11 -127
rect -80 -139 -68 -135
rect -97 -228 -93 -151
rect -80 -159 -76 -139
rect -48 -147 -40 -143
rect -37 -143 -34 -131
rect -37 -147 -30 -143
rect -43 -151 -40 -147
rect -43 -155 -30 -151
rect -15 -159 -11 -131
rect -8 -131 -4 -111
rect 8 -121 12 -101
rect 15 -109 19 -65
rect 22 -73 29 -69
rect 82 -71 85 -69
rect 78 -73 85 -71
rect 22 -101 25 -73
rect 78 -77 82 -73
rect 69 -81 82 -77
rect 69 -97 75 -93
rect 22 -105 29 -101
rect 71 -109 75 -97
rect 78 -101 82 -81
rect 111 -85 115 -49
rect 105 -89 111 -85
rect 78 -105 85 -101
rect 15 -113 75 -109
rect 15 -125 19 -113
rect 48 -121 90 -117
rect 111 -125 115 -89
rect 15 -129 28 -125
rect 100 -129 115 -125
rect 15 -145 19 -129
rect 48 -141 95 -137
rect 15 -149 28 -145
rect 111 -145 115 -129
rect 15 -154 19 -149
rect 60 -154 64 -148
rect 105 -149 115 -145
rect 129 -149 132 -106
rect 15 -158 28 -154
rect 60 -158 87 -154
rect -80 -163 -68 -159
rect -20 -163 -15 -159
rect 0 -162 8 -158
rect 0 -163 4 -162
rect -80 -176 -76 -163
rect -48 -169 -39 -168
rect -34 -169 -30 -168
rect -48 -172 -30 -169
rect -80 -180 -68 -176
rect -15 -176 -11 -163
rect -80 -184 -76 -180
rect -39 -184 -35 -179
rect -20 -180 -11 -176
rect -80 -188 -68 -184
rect -44 -187 -30 -184
rect -80 -200 -76 -188
rect -44 -192 -41 -187
rect -48 -196 -41 -192
rect -80 -204 -68 -200
rect -15 -200 -11 -180
rect -87 -228 -83 -216
rect -97 -232 -87 -228
rect -80 -216 -76 -204
rect -38 -208 -34 -203
rect -20 -204 -11 -200
rect -15 -208 -11 -204
rect -48 -212 -34 -208
rect -20 -212 -11 -208
rect -80 -220 -68 -216
rect -97 -309 -93 -232
rect -80 -240 -76 -220
rect -48 -228 -40 -224
rect -37 -224 -34 -212
rect -37 -228 -30 -224
rect -43 -232 -40 -228
rect -43 -236 -30 -232
rect -15 -240 -11 -212
rect -8 -212 -4 -192
rect 0 -232 4 -168
rect 8 -184 12 -170
rect 8 -202 12 -188
rect 8 -224 12 -207
rect 15 -170 19 -158
rect 73 -162 77 -158
rect 48 -166 77 -162
rect 111 -170 115 -149
rect 15 -174 28 -170
rect 107 -174 115 -170
rect 15 -180 19 -174
rect 111 -180 115 -174
rect 15 -184 28 -180
rect 100 -184 115 -180
rect 15 -196 19 -184
rect 48 -192 90 -188
rect 15 -200 25 -196
rect 0 -236 8 -232
rect -80 -244 -68 -240
rect -20 -244 -15 -240
rect -80 -257 -76 -244
rect -48 -253 -30 -249
rect -80 -261 -68 -257
rect -15 -257 -11 -244
rect -80 -265 -76 -261
rect -39 -265 -35 -260
rect -20 -261 -11 -257
rect 8 -256 12 -236
rect 15 -244 19 -200
rect 22 -208 29 -204
rect 82 -206 85 -204
rect 78 -208 85 -206
rect 22 -236 25 -208
rect 78 -212 82 -208
rect 69 -216 82 -212
rect 69 -232 75 -228
rect 22 -240 29 -236
rect 71 -244 75 -232
rect 78 -236 82 -216
rect 111 -220 115 -184
rect 105 -224 111 -220
rect 78 -240 85 -236
rect 15 -248 75 -244
rect 15 -260 19 -248
rect 48 -256 90 -252
rect 111 -260 115 -224
rect 127 -220 133 -217
rect -80 -269 -68 -265
rect -44 -268 -30 -265
rect -80 -281 -76 -269
rect -44 -273 -41 -268
rect -48 -277 -41 -273
rect -80 -285 -68 -281
rect -15 -281 -11 -261
rect 15 -264 28 -260
rect 100 -264 115 -260
rect -87 -309 -83 -297
rect -97 -313 -87 -309
rect -80 -297 -76 -285
rect -38 -289 -34 -284
rect -20 -285 -11 -281
rect -15 -289 -11 -285
rect -48 -293 -34 -289
rect -20 -293 -11 -289
rect -80 -301 -68 -297
rect -97 -389 -93 -313
rect -80 -321 -76 -301
rect -48 -309 -40 -305
rect -37 -305 -34 -293
rect -37 -309 -30 -305
rect -43 -313 -40 -309
rect -43 -317 -30 -313
rect -15 -321 -11 -293
rect -8 -293 -4 -273
rect 15 -277 19 -264
rect 48 -273 95 -269
rect 15 -281 28 -277
rect 111 -277 115 -264
rect 15 -286 19 -281
rect 60 -286 64 -280
rect 105 -281 115 -277
rect 127 -281 130 -220
rect 15 -290 28 -286
rect 60 -290 87 -286
rect 0 -294 8 -290
rect -80 -325 -68 -321
rect -20 -325 -15 -321
rect 0 -324 4 -294
rect -80 -337 -76 -325
rect -48 -330 -39 -329
rect -34 -330 -30 -329
rect -48 -333 -30 -330
rect -80 -341 -68 -337
rect -15 -337 -11 -325
rect -80 -345 -76 -341
rect -39 -345 -35 -340
rect -20 -341 -11 -337
rect -80 -349 -68 -345
rect -44 -348 -30 -345
rect -80 -361 -76 -349
rect -44 -353 -41 -348
rect -48 -357 -41 -353
rect -80 -365 -68 -361
rect -15 -361 -11 -341
rect -87 -389 -83 -377
rect -97 -393 -87 -389
rect -80 -377 -76 -365
rect -38 -369 -34 -364
rect -20 -365 -11 -361
rect -15 -369 -11 -365
rect -48 -373 -34 -369
rect -20 -373 -11 -369
rect -80 -381 -68 -377
rect -97 -470 -93 -393
rect -80 -401 -76 -381
rect -48 -389 -40 -385
rect -37 -385 -34 -373
rect -37 -389 -30 -385
rect -43 -393 -40 -389
rect -43 -397 -30 -393
rect -15 -401 -11 -373
rect -8 -373 -4 -353
rect 0 -364 4 -329
rect 8 -316 12 -302
rect 8 -341 12 -320
rect 8 -356 12 -346
rect 15 -302 19 -290
rect 73 -294 77 -290
rect 48 -298 77 -294
rect 111 -302 115 -281
rect 15 -306 28 -302
rect 107 -306 115 -302
rect 15 -312 19 -306
rect 111 -312 115 -306
rect 15 -316 28 -312
rect 100 -316 115 -312
rect 15 -328 19 -316
rect 48 -324 90 -320
rect 15 -332 25 -328
rect 0 -368 8 -364
rect 8 -388 12 -368
rect 15 -376 19 -332
rect 22 -340 29 -336
rect 82 -338 85 -336
rect 78 -340 85 -338
rect 22 -368 25 -340
rect 78 -344 82 -340
rect 69 -348 82 -344
rect 69 -364 75 -360
rect 22 -372 29 -368
rect 71 -376 75 -364
rect 78 -368 82 -348
rect 111 -352 115 -316
rect 105 -356 111 -352
rect 78 -372 85 -368
rect 15 -380 75 -376
rect 15 -392 19 -380
rect 48 -388 90 -384
rect 111 -392 115 -356
rect -80 -405 -68 -401
rect -20 -405 -15 -401
rect -80 -418 -76 -405
rect -48 -414 -30 -410
rect -80 -422 -68 -418
rect -15 -418 -11 -405
rect -80 -426 -76 -422
rect -39 -426 -35 -421
rect -20 -422 -11 -418
rect -80 -430 -68 -426
rect -44 -429 -30 -426
rect -80 -442 -76 -430
rect -44 -434 -41 -429
rect -48 -438 -41 -434
rect -80 -446 -68 -442
rect -15 -442 -11 -422
rect 15 -396 28 -392
rect 100 -396 115 -392
rect 15 -411 19 -396
rect 48 -407 95 -403
rect 15 -415 28 -411
rect 111 -411 115 -396
rect 15 -420 19 -415
rect 60 -420 64 -414
rect 105 -415 115 -411
rect 15 -424 28 -420
rect 60 -424 87 -420
rect 0 -428 8 -424
rect -87 -470 -83 -458
rect -97 -474 -87 -470
rect -80 -458 -76 -446
rect -38 -450 -34 -445
rect -20 -446 -11 -442
rect -15 -450 -11 -446
rect -48 -454 -34 -450
rect -20 -454 -11 -450
rect -80 -462 -68 -458
rect -97 -551 -93 -474
rect -80 -482 -76 -462
rect -48 -470 -40 -466
rect -37 -466 -34 -454
rect -37 -470 -30 -466
rect -43 -474 -40 -470
rect -43 -478 -30 -474
rect -15 -482 -11 -454
rect -8 -454 -4 -434
rect -80 -486 -68 -482
rect -20 -486 -15 -482
rect -80 -499 -76 -486
rect -48 -492 -40 -491
rect -35 -492 -30 -491
rect -48 -495 -30 -492
rect -80 -503 -68 -499
rect -15 -499 -11 -487
rect -80 -507 -76 -503
rect -39 -507 -35 -502
rect -20 -503 -11 -499
rect -80 -511 -68 -507
rect -44 -510 -30 -507
rect -80 -523 -76 -511
rect -44 -515 -41 -510
rect -48 -519 -41 -515
rect -80 -527 -68 -523
rect -15 -523 -11 -503
rect -8 -500 -4 -479
rect 0 -487 4 -428
rect 8 -450 12 -436
rect 8 -474 12 -454
rect 0 -498 4 -492
rect 8 -490 12 -479
rect 15 -436 19 -424
rect 73 -428 77 -424
rect 48 -432 77 -428
rect 111 -436 115 -415
rect 15 -440 28 -436
rect 107 -440 115 -436
rect 15 -446 19 -440
rect 111 -446 115 -440
rect 15 -450 28 -446
rect 100 -450 115 -446
rect 15 -462 19 -450
rect 48 -458 90 -454
rect 15 -466 25 -462
rect 0 -502 8 -498
rect -87 -551 -83 -539
rect -97 -555 -87 -551
rect -80 -539 -76 -527
rect -38 -531 -34 -526
rect -20 -527 -11 -523
rect -15 -531 -11 -527
rect -48 -535 -34 -531
rect -20 -535 -11 -531
rect -80 -543 -68 -539
rect -97 -632 -93 -555
rect -80 -563 -76 -543
rect -48 -551 -40 -547
rect -37 -547 -34 -535
rect -37 -551 -30 -547
rect -43 -555 -40 -551
rect -43 -559 -30 -555
rect -15 -563 -11 -535
rect -8 -535 -4 -515
rect 8 -522 12 -502
rect 15 -510 19 -466
rect 22 -474 29 -470
rect 82 -472 85 -470
rect 78 -474 85 -472
rect 22 -502 25 -474
rect 78 -478 82 -474
rect 69 -482 82 -478
rect 69 -498 75 -494
rect 22 -506 29 -502
rect 71 -510 75 -498
rect 78 -502 82 -482
rect 111 -486 115 -450
rect 105 -490 111 -486
rect 78 -506 85 -502
rect 15 -514 75 -510
rect 15 -526 19 -514
rect 48 -522 90 -518
rect 111 -526 115 -490
rect 128 -490 131 -446
rect 15 -530 28 -526
rect 100 -530 115 -526
rect 15 -535 19 -530
rect -80 -567 -68 -563
rect -20 -567 -15 -563
rect -80 -580 -76 -567
rect -48 -576 -30 -572
rect -80 -584 -68 -580
rect -15 -580 -11 -567
rect -80 -588 -76 -584
rect -39 -588 -35 -583
rect -20 -584 -11 -580
rect -15 -585 -11 -584
rect 111 -585 115 -530
rect 128 -531 131 -496
rect 128 -564 131 -537
rect -80 -592 -68 -588
rect -44 -591 -30 -588
rect -80 -604 -76 -592
rect -44 -596 -41 -591
rect -15 -589 115 -585
rect -48 -600 -41 -596
rect -80 -608 -68 -604
rect -15 -604 -11 -589
rect -87 -632 -83 -620
rect -97 -636 -87 -632
rect -80 -620 -76 -608
rect -38 -612 -34 -607
rect -20 -608 -11 -604
rect -15 -612 -11 -608
rect -48 -616 -34 -612
rect -20 -616 -11 -612
rect -80 -624 -68 -620
rect -97 -653 -93 -636
rect -80 -644 -76 -624
rect -48 -632 -40 -628
rect -37 -628 -34 -616
rect -37 -632 -30 -628
rect -43 -636 -40 -632
rect -43 -640 -30 -636
rect -15 -644 -11 -616
rect -8 -616 -4 -596
rect 111 -609 115 -589
rect 128 -590 131 -570
rect 135 -582 138 -273
rect 142 -307 145 -232
rect 142 -342 145 -312
rect 142 -367 145 -347
rect 149 -358 152 -136
rect 156 -201 159 -180
rect 163 -192 166 -2
rect 170 -59 173 -45
rect 170 -84 173 -64
rect 177 -75 180 130
rect 184 -8 187 87
rect 191 0 194 130
rect 209 41 213 146
rect 286 130 290 141
rect 310 137 314 141
rect 302 134 314 137
rect 302 132 305 134
rect 276 126 290 130
rect 297 128 305 132
rect 326 131 330 141
rect 342 136 346 141
rect 342 133 354 136
rect 286 123 290 126
rect 302 123 305 128
rect 321 130 330 131
rect 321 127 346 130
rect 342 123 346 127
rect 350 123 354 133
rect 220 49 223 113
rect 294 108 298 113
rect 318 108 322 113
rect 326 108 330 113
rect 358 108 362 113
rect 276 104 358 108
rect 310 97 330 101
rect 372 65 376 169
rect 372 61 508 65
rect 209 37 495 41
rect 209 12 213 37
rect 209 8 218 12
rect 209 4 213 8
rect 330 4 334 26
rect 209 0 221 4
rect 277 0 330 4
rect 191 -4 202 0
rect 184 -50 187 -13
rect 191 -43 194 -4
rect 209 -12 213 0
rect 241 -8 253 -4
rect 249 -12 253 -8
rect 209 -16 221 -12
rect 249 -16 257 -12
rect 261 -16 321 -12
rect 209 -31 213 -16
rect 209 -35 219 -31
rect 191 -47 202 -43
rect 209 -47 213 -35
rect 330 -39 334 0
rect 348 -4 352 15
rect 355 8 359 37
rect 355 4 364 8
rect 355 0 359 4
rect 472 0 476 27
rect 355 -4 367 0
rect 421 -4 472 0
rect 355 -16 359 -4
rect 387 -12 394 -8
rect 355 -20 367 -16
rect 391 -20 394 -12
rect 398 -20 401 -16
rect 241 -43 253 -39
rect 287 -43 334 -39
rect 170 -135 173 -89
rect 170 -167 173 -140
rect 177 -158 180 -80
rect 184 -126 187 -55
rect 191 -119 194 -47
rect 209 -51 221 -47
rect 209 -63 213 -51
rect 249 -55 253 -43
rect 241 -59 253 -55
rect 249 -63 253 -59
rect 209 -67 221 -63
rect 249 -67 257 -63
rect 261 -67 321 -63
rect 209 -72 213 -67
rect 330 -72 334 -43
rect 348 -67 352 -26
rect 355 -55 359 -20
rect 391 -23 401 -20
rect 397 -28 401 -23
rect 355 -59 364 -55
rect 355 -71 359 -59
rect 472 -63 476 -4
rect 491 23 495 37
rect 504 34 508 61
rect 504 30 600 34
rect 491 19 626 23
rect 491 -13 495 19
rect 587 -13 591 -7
rect 491 -17 504 -13
rect 576 -17 591 -13
rect 484 -35 488 -21
rect 484 -57 488 -40
rect 491 -29 495 -17
rect 524 -25 566 -21
rect 491 -33 501 -29
rect 387 -67 400 -63
rect 433 -67 472 -63
rect 209 -76 221 -72
rect 277 -76 334 -72
rect 355 -75 367 -71
rect 209 -88 213 -76
rect 241 -84 253 -80
rect 249 -88 253 -84
rect 209 -92 221 -88
rect 249 -92 257 -88
rect 261 -92 321 -88
rect 209 -107 213 -92
rect 209 -111 218 -107
rect 209 -115 213 -111
rect 330 -115 334 -76
rect 355 -87 359 -75
rect 396 -79 400 -67
rect 387 -83 400 -79
rect 396 -87 400 -83
rect 355 -91 367 -87
rect 396 -91 403 -87
rect 209 -119 221 -115
rect 296 -119 334 -115
rect 191 -123 202 -119
rect 156 -260 159 -206
rect 156 -300 159 -265
rect 156 -333 159 -305
rect 163 -324 166 -197
rect 170 -251 173 -172
rect 170 -292 173 -256
rect 142 -433 145 -372
rect 142 -482 145 -438
rect 142 -522 145 -487
rect 142 -557 145 -528
rect 149 -549 152 -363
rect 156 -425 159 -338
rect 156 -474 159 -430
rect 156 -516 159 -479
rect 163 -508 166 -329
rect 170 -417 173 -297
rect 170 -467 173 -422
rect 177 -459 180 -163
rect 184 -243 187 -131
rect 191 -235 194 -123
rect 209 -131 213 -119
rect 241 -127 253 -123
rect 209 -135 221 -131
rect 209 -147 213 -135
rect 249 -139 253 -127
rect 241 -143 253 -139
rect 249 -147 253 -143
rect 209 -151 221 -147
rect 249 -151 256 -147
rect 260 -151 321 -147
rect 209 -164 213 -151
rect 330 -156 334 -119
rect 241 -160 253 -156
rect 286 -160 334 -156
rect 209 -168 221 -164
rect 209 -180 213 -168
rect 249 -172 253 -160
rect 241 -176 253 -172
rect 249 -180 253 -176
rect 209 -184 221 -180
rect 249 -184 256 -180
rect 260 -184 321 -180
rect 209 -189 213 -184
rect 330 -189 334 -160
rect 347 -164 351 -106
rect 355 -152 359 -91
rect 396 -94 400 -91
rect 355 -156 364 -152
rect 355 -160 359 -156
rect 472 -160 476 -67
rect 484 -78 488 -69
rect 484 -89 488 -83
rect 491 -77 495 -33
rect 498 -41 505 -37
rect 558 -39 561 -37
rect 554 -41 561 -39
rect 498 -69 501 -41
rect 554 -45 558 -41
rect 545 -49 558 -45
rect 545 -65 551 -61
rect 498 -73 505 -69
rect 547 -77 551 -65
rect 554 -69 558 -49
rect 587 -53 591 -17
rect 602 -45 606 6
rect 622 7 626 19
rect 654 11 672 15
rect 622 3 634 7
rect 687 7 691 19
rect 622 -1 626 3
rect 663 -1 667 4
rect 682 3 691 7
rect 622 -5 634 -1
rect 658 -4 672 -1
rect 622 -17 626 -5
rect 658 -9 661 -4
rect 654 -13 661 -9
rect 622 -21 634 -17
rect 687 -17 691 3
rect 615 -45 619 -33
rect 602 -49 615 -45
rect 622 -33 626 -21
rect 664 -25 668 -20
rect 682 -21 691 -17
rect 687 -25 691 -21
rect 654 -29 668 -25
rect 682 -29 691 -25
rect 622 -37 634 -33
rect 581 -57 587 -53
rect 554 -73 561 -69
rect 491 -81 551 -77
rect 491 -93 495 -81
rect 524 -89 566 -85
rect 587 -93 591 -57
rect 491 -97 504 -93
rect 576 -97 591 -93
rect 491 -103 495 -97
rect 587 -103 591 -97
rect 491 -107 504 -103
rect 576 -107 591 -103
rect 484 -126 488 -111
rect 484 -147 488 -131
rect 491 -119 495 -107
rect 524 -115 566 -111
rect 491 -123 501 -119
rect 355 -164 367 -160
rect 432 -164 472 -160
rect 355 -176 359 -164
rect 387 -172 399 -168
rect 355 -180 367 -176
rect 209 -193 221 -189
rect 276 -193 334 -189
rect 209 -205 213 -193
rect 241 -201 253 -197
rect 249 -205 253 -201
rect 209 -209 221 -205
rect 249 -209 256 -205
rect 260 -209 321 -205
rect 209 -224 213 -209
rect 209 -228 218 -224
rect 191 -239 202 -235
rect 184 -284 187 -248
rect 184 -410 187 -289
rect 191 -402 194 -239
rect 209 -240 213 -228
rect 330 -232 334 -193
rect 355 -192 359 -180
rect 395 -184 399 -172
rect 387 -188 399 -184
rect 395 -192 399 -188
rect 355 -196 367 -192
rect 395 -196 402 -192
rect 241 -236 253 -232
rect 306 -236 334 -232
rect 209 -244 221 -240
rect 209 -256 213 -244
rect 249 -248 253 -236
rect 241 -252 253 -248
rect 209 -260 221 -256
rect 209 -272 213 -260
rect 249 -264 253 -252
rect 241 -268 253 -264
rect 249 -272 253 -268
rect 209 -276 221 -272
rect 249 -276 256 -272
rect 260 -276 321 -272
rect 209 -281 213 -276
rect 330 -281 334 -236
rect 209 -285 221 -281
rect 296 -285 334 -281
rect 209 -297 213 -285
rect 241 -293 253 -289
rect 209 -301 221 -297
rect 209 -313 213 -301
rect 249 -305 253 -293
rect 241 -309 253 -305
rect 249 -313 253 -309
rect 209 -317 221 -313
rect 249 -317 256 -313
rect 260 -317 321 -313
rect 209 -330 213 -317
rect 330 -322 334 -285
rect 340 -314 344 -277
rect 347 -306 351 -221
rect 355 -294 359 -196
rect 395 -199 399 -196
rect 355 -298 364 -294
rect 355 -310 359 -298
rect 472 -302 476 -164
rect 484 -167 488 -159
rect 484 -179 488 -172
rect 491 -167 495 -123
rect 498 -131 505 -127
rect 558 -129 561 -127
rect 554 -131 561 -129
rect 498 -159 501 -131
rect 554 -135 558 -131
rect 545 -139 558 -135
rect 545 -155 551 -151
rect 498 -163 505 -159
rect 547 -167 551 -155
rect 554 -159 558 -139
rect 587 -143 591 -107
rect 602 -126 606 -49
rect 622 -57 626 -37
rect 654 -45 662 -41
rect 665 -41 668 -29
rect 665 -45 672 -41
rect 659 -49 662 -45
rect 659 -53 672 -49
rect 687 -57 691 -29
rect 694 -29 698 -9
rect 622 -61 634 -57
rect 682 -61 687 -57
rect 622 -74 626 -61
rect 654 -70 672 -66
rect 622 -78 634 -74
rect 687 -74 691 -61
rect 622 -82 626 -78
rect 663 -82 667 -77
rect 682 -78 691 -74
rect 622 -86 634 -82
rect 658 -85 672 -82
rect 622 -98 626 -86
rect 658 -90 661 -85
rect 654 -94 661 -90
rect 622 -102 634 -98
rect 687 -98 691 -78
rect 615 -126 619 -114
rect 602 -130 615 -126
rect 622 -114 626 -102
rect 664 -106 668 -101
rect 682 -102 691 -98
rect 687 -106 691 -102
rect 654 -110 668 -106
rect 682 -110 691 -106
rect 622 -118 634 -114
rect 581 -147 587 -143
rect 554 -163 561 -159
rect 491 -171 551 -167
rect 491 -183 495 -171
rect 524 -179 566 -175
rect 587 -183 591 -147
rect 491 -187 504 -183
rect 576 -187 591 -183
rect 491 -192 495 -187
rect 587 -192 591 -187
rect 491 -196 504 -192
rect 576 -196 591 -192
rect 484 -218 488 -200
rect 484 -236 488 -223
rect 491 -208 495 -196
rect 524 -204 566 -200
rect 491 -212 501 -208
rect 484 -258 488 -248
rect 484 -268 488 -263
rect 491 -256 495 -212
rect 498 -220 505 -216
rect 558 -218 561 -216
rect 554 -220 561 -218
rect 498 -248 501 -220
rect 554 -224 558 -220
rect 545 -228 558 -224
rect 545 -244 551 -240
rect 498 -252 505 -248
rect 547 -256 551 -244
rect 554 -248 558 -228
rect 587 -232 591 -196
rect 602 -207 606 -130
rect 622 -138 626 -118
rect 654 -126 662 -122
rect 665 -122 668 -110
rect 665 -126 672 -122
rect 659 -130 662 -126
rect 659 -134 672 -130
rect 687 -138 691 -110
rect 694 -110 698 -90
rect 622 -142 634 -138
rect 682 -142 687 -138
rect 622 -155 626 -142
rect 654 -151 672 -147
rect 622 -159 634 -155
rect 687 -155 691 -143
rect 622 -163 626 -159
rect 663 -163 667 -158
rect 682 -159 691 -155
rect 622 -167 634 -163
rect 658 -166 672 -163
rect 622 -179 626 -167
rect 658 -171 661 -166
rect 654 -175 661 -171
rect 622 -183 634 -179
rect 687 -179 691 -159
rect 615 -207 619 -195
rect 602 -211 615 -207
rect 622 -195 626 -183
rect 664 -187 668 -182
rect 682 -183 691 -179
rect 687 -187 691 -183
rect 654 -191 668 -187
rect 682 -191 691 -187
rect 622 -199 634 -195
rect 581 -236 587 -232
rect 554 -252 561 -248
rect 491 -260 551 -256
rect 491 -272 495 -260
rect 524 -268 566 -264
rect 587 -272 591 -236
rect 491 -276 504 -272
rect 576 -276 591 -272
rect 491 -280 495 -276
rect 587 -280 591 -276
rect 491 -284 504 -280
rect 576 -284 591 -280
rect 388 -306 399 -302
rect 442 -306 472 -302
rect 355 -314 368 -310
rect 340 -318 347 -314
rect 241 -326 253 -322
rect 286 -326 334 -322
rect 355 -326 359 -314
rect 395 -318 399 -306
rect 388 -322 399 -318
rect 209 -334 221 -330
rect 209 -346 213 -334
rect 249 -338 253 -326
rect 241 -342 253 -338
rect 249 -346 253 -342
rect 209 -350 221 -346
rect 249 -350 256 -346
rect 260 -350 321 -346
rect 209 -355 213 -350
rect 330 -355 334 -326
rect 355 -330 368 -326
rect 355 -342 359 -330
rect 395 -334 399 -322
rect 388 -338 399 -334
rect 395 -342 399 -338
rect 355 -346 368 -342
rect 395 -346 402 -342
rect 209 -359 221 -355
rect 276 -359 334 -355
rect 209 -371 213 -359
rect 241 -367 253 -363
rect 249 -371 253 -367
rect 209 -375 221 -371
rect 249 -375 256 -371
rect 260 -375 321 -371
rect 209 -390 213 -375
rect 209 -394 218 -390
rect 209 -398 213 -394
rect 330 -398 334 -359
rect 209 -402 221 -398
rect 316 -402 334 -398
rect 191 -406 202 -402
rect 184 -414 202 -410
rect 209 -414 213 -402
rect 241 -410 253 -406
rect 209 -418 221 -414
rect 193 -430 202 -426
rect 209 -430 213 -418
rect 249 -422 253 -410
rect 241 -426 253 -422
rect 209 -434 221 -430
rect 209 -446 213 -434
rect 249 -438 253 -426
rect 241 -442 253 -438
rect 249 -446 253 -442
rect 209 -450 221 -446
rect 249 -450 256 -446
rect 260 -450 321 -446
rect 177 -463 202 -459
rect 209 -463 213 -450
rect 330 -455 334 -402
rect 241 -459 253 -455
rect 306 -459 334 -455
rect 209 -467 221 -463
rect 170 -471 202 -467
rect 182 -479 202 -475
rect 209 -479 213 -467
rect 249 -471 253 -459
rect 241 -475 253 -471
rect 209 -483 221 -479
rect 209 -495 213 -483
rect 249 -487 253 -475
rect 241 -491 253 -487
rect 249 -495 253 -491
rect 209 -499 221 -495
rect 249 -499 256 -495
rect 260 -499 321 -495
rect 209 -504 213 -499
rect 330 -504 334 -459
rect 209 -508 221 -504
rect 296 -508 334 -504
rect 163 -512 202 -508
rect 156 -520 202 -516
rect 209 -520 213 -508
rect 241 -516 253 -512
rect 209 -524 221 -520
rect 209 -536 213 -524
rect 249 -528 253 -516
rect 241 -532 253 -528
rect 249 -536 253 -532
rect 209 -540 221 -536
rect 249 -540 256 -536
rect 260 -540 321 -536
rect 149 -553 202 -549
rect 209 -553 213 -540
rect 330 -545 334 -508
rect 340 -520 344 -451
rect 347 -512 351 -386
rect 355 -500 359 -346
rect 395 -351 399 -346
rect 397 -499 462 -496
rect 355 -504 365 -500
rect 355 -508 359 -504
rect 355 -512 368 -508
rect 340 -523 347 -520
rect 355 -524 359 -512
rect 397 -516 401 -499
rect 472 -508 476 -306
rect 484 -324 488 -293
rect 491 -296 495 -284
rect 524 -292 566 -288
rect 491 -300 501 -296
rect 484 -342 488 -336
rect 484 -356 488 -347
rect 491 -344 495 -300
rect 498 -308 505 -304
rect 558 -306 561 -304
rect 554 -308 561 -306
rect 498 -336 501 -308
rect 554 -312 558 -308
rect 545 -316 558 -312
rect 545 -332 551 -328
rect 498 -340 505 -336
rect 547 -344 551 -332
rect 554 -336 558 -316
rect 587 -320 591 -284
rect 602 -288 606 -211
rect 622 -219 626 -199
rect 654 -207 662 -203
rect 665 -203 668 -191
rect 665 -207 672 -203
rect 659 -211 662 -207
rect 659 -215 672 -211
rect 687 -219 691 -191
rect 694 -191 698 -171
rect 622 -223 634 -219
rect 682 -223 687 -219
rect 622 -236 626 -223
rect 654 -232 672 -228
rect 622 -240 634 -236
rect 687 -236 691 -223
rect 622 -244 626 -240
rect 663 -244 667 -239
rect 682 -240 691 -236
rect 622 -248 634 -244
rect 658 -247 672 -244
rect 622 -260 626 -248
rect 658 -252 661 -247
rect 654 -256 661 -252
rect 622 -264 634 -260
rect 687 -260 691 -240
rect 615 -288 619 -276
rect 602 -292 615 -288
rect 622 -276 626 -264
rect 664 -268 668 -263
rect 682 -264 691 -260
rect 687 -268 691 -264
rect 654 -272 668 -268
rect 682 -272 691 -268
rect 622 -280 634 -276
rect 581 -324 587 -320
rect 554 -340 561 -336
rect 491 -348 551 -344
rect 491 -360 495 -348
rect 524 -356 566 -352
rect 587 -360 591 -324
rect 491 -364 504 -360
rect 576 -364 591 -360
rect 491 -369 495 -364
rect 587 -369 591 -364
rect 491 -373 504 -369
rect 576 -373 591 -369
rect 484 -400 488 -377
rect 484 -413 488 -405
rect 491 -385 495 -373
rect 524 -381 566 -377
rect 491 -389 501 -385
rect 484 -430 488 -425
rect 484 -445 488 -435
rect 491 -433 495 -389
rect 498 -397 505 -393
rect 558 -395 561 -393
rect 554 -397 561 -395
rect 498 -425 501 -397
rect 554 -401 558 -397
rect 545 -405 558 -401
rect 545 -421 551 -417
rect 498 -429 505 -425
rect 547 -433 551 -421
rect 554 -425 558 -405
rect 587 -409 591 -373
rect 602 -369 606 -292
rect 622 -300 626 -280
rect 654 -288 662 -284
rect 665 -284 668 -272
rect 665 -288 672 -284
rect 659 -292 662 -288
rect 659 -296 672 -292
rect 687 -300 691 -272
rect 694 -272 698 -252
rect 622 -304 634 -300
rect 682 -304 687 -300
rect 622 -317 626 -304
rect 654 -313 672 -309
rect 622 -321 634 -317
rect 687 -317 691 -305
rect 622 -325 626 -321
rect 663 -325 667 -320
rect 682 -321 691 -317
rect 622 -329 634 -325
rect 658 -328 672 -325
rect 622 -341 626 -329
rect 658 -333 661 -328
rect 654 -337 661 -333
rect 622 -345 634 -341
rect 687 -341 691 -321
rect 615 -369 619 -357
rect 602 -373 615 -369
rect 622 -357 626 -345
rect 664 -349 668 -344
rect 682 -345 691 -341
rect 687 -349 691 -345
rect 654 -353 668 -349
rect 682 -353 691 -349
rect 622 -361 634 -357
rect 581 -413 587 -409
rect 554 -429 561 -425
rect 491 -437 551 -433
rect 491 -449 495 -437
rect 524 -445 566 -441
rect 587 -449 591 -413
rect 491 -453 504 -449
rect 576 -453 591 -449
rect 491 -459 495 -453
rect 587 -470 591 -453
rect 602 -450 606 -373
rect 622 -381 626 -361
rect 654 -369 662 -365
rect 665 -365 668 -353
rect 665 -369 672 -365
rect 659 -373 662 -369
rect 659 -377 672 -373
rect 687 -381 691 -353
rect 694 -353 698 -333
rect 622 -385 634 -381
rect 682 -385 687 -381
rect 622 -398 626 -385
rect 654 -394 672 -390
rect 622 -402 634 -398
rect 687 -398 691 -385
rect 622 -406 626 -402
rect 663 -406 667 -401
rect 682 -402 691 -398
rect 622 -410 634 -406
rect 658 -409 672 -406
rect 622 -422 626 -410
rect 658 -414 661 -409
rect 654 -418 661 -414
rect 622 -426 634 -422
rect 687 -422 691 -402
rect 615 -450 619 -438
rect 602 -454 615 -450
rect 622 -438 626 -426
rect 664 -430 668 -425
rect 682 -426 691 -422
rect 687 -430 691 -426
rect 654 -434 668 -430
rect 682 -434 691 -430
rect 622 -442 634 -438
rect 622 -462 626 -442
rect 654 -450 662 -446
rect 665 -446 668 -434
rect 665 -450 672 -446
rect 659 -454 662 -450
rect 659 -458 672 -454
rect 687 -462 691 -434
rect 694 -434 698 -414
rect 622 -466 634 -462
rect 682 -466 687 -462
rect 622 -472 626 -466
rect 587 -482 591 -474
rect 687 -482 691 -466
rect 587 -486 691 -482
rect 465 -512 472 -508
rect 388 -520 401 -516
rect 355 -528 368 -524
rect 342 -532 347 -528
rect 355 -540 359 -528
rect 397 -532 401 -520
rect 388 -536 401 -532
rect 355 -544 368 -540
rect 241 -549 253 -545
rect 286 -549 334 -545
rect 344 -548 347 -544
rect 209 -557 221 -553
rect 142 -561 202 -557
rect 209 -569 213 -557
rect 249 -561 253 -549
rect 241 -565 253 -561
rect 249 -569 253 -565
rect 209 -573 221 -569
rect 249 -573 256 -569
rect 260 -573 321 -569
rect 209 -578 213 -573
rect 330 -578 334 -549
rect 355 -556 359 -544
rect 397 -548 401 -536
rect 388 -552 401 -548
rect 397 -556 401 -552
rect 355 -560 368 -556
rect 397 -560 405 -556
rect 355 -568 359 -560
rect 209 -582 221 -578
rect 276 -582 334 -578
rect 135 -586 202 -582
rect 128 -594 202 -590
rect 209 -594 213 -582
rect 241 -590 253 -586
rect 249 -594 253 -590
rect 209 -598 221 -594
rect 249 -598 256 -594
rect 260 -598 321 -594
rect 209 -604 213 -598
rect 330 -609 334 -582
rect 472 -609 476 -512
rect 479 -507 483 -506
rect 587 -507 591 -486
rect 479 -511 591 -507
rect 479 -609 483 -511
rect 111 -613 483 -609
rect -80 -648 -68 -644
rect -20 -648 -15 -644
rect -80 -654 -76 -648
<< m2contact >>
rect -38 74 -33 79
rect 59 130 65 135
rect 176 130 181 135
rect 190 130 195 135
rect 73 113 78 118
rect 7 74 12 79
rect 94 74 99 79
rect 77 61 82 66
rect 118 59 123 64
rect 94 11 99 16
rect 118 42 123 47
rect -39 -7 -34 -2
rect 0 -6 5 -1
rect 59 -2 65 3
rect 162 -2 167 3
rect 73 -19 78 -14
rect -38 -87 -33 -82
rect 7 -87 12 -82
rect 94 -58 99 -53
rect 77 -71 82 -66
rect 118 -73 123 -68
rect 94 -121 99 -116
rect 118 -90 123 -85
rect 128 -106 133 -101
rect 59 -137 65 -132
rect 148 -136 153 -131
rect 73 -154 78 -149
rect -39 -169 -34 -164
rect -1 -168 4 -163
rect 7 -207 12 -202
rect 128 -154 133 -149
rect 94 -193 99 -188
rect -38 -249 -33 -244
rect 77 -206 82 -201
rect 118 -208 123 -203
rect 94 -256 99 -251
rect 118 -225 123 -220
rect 59 -269 65 -264
rect 133 -221 138 -216
rect 141 -232 146 -227
rect 134 -273 139 -268
rect 73 -286 78 -281
rect -39 -330 -34 -325
rect -1 -329 4 -324
rect 7 -346 12 -341
rect 126 -286 131 -281
rect 94 -325 99 -320
rect 77 -338 82 -333
rect 118 -340 123 -335
rect 94 -388 99 -383
rect 118 -357 123 -352
rect -38 -410 -33 -405
rect 59 -403 65 -398
rect 73 -420 78 -415
rect -40 -492 -35 -487
rect -8 -479 -3 -474
rect 7 -479 12 -474
rect -1 -492 4 -487
rect 127 -446 132 -441
rect 94 -459 99 -454
rect -8 -505 -3 -500
rect 77 -472 82 -467
rect 118 -474 123 -469
rect 94 -522 99 -517
rect 118 -491 123 -486
rect 127 -496 132 -490
rect -38 -572 -33 -567
rect 127 -537 132 -531
rect 127 -570 132 -564
rect 141 -312 146 -307
rect 141 -347 146 -342
rect 155 -180 160 -175
rect 169 -45 174 -40
rect 169 -64 174 -59
rect 183 87 188 92
rect 219 113 224 118
rect 219 44 224 49
rect 347 15 352 20
rect 183 -13 188 -8
rect 197 -13 202 -8
rect 321 -17 326 -12
rect 343 -17 348 -12
rect 347 -26 352 -21
rect 183 -55 188 -50
rect 176 -80 181 -75
rect 169 -89 174 -84
rect 169 -140 174 -135
rect 197 -55 202 -50
rect 197 -64 202 -59
rect 321 -68 326 -63
rect 396 -33 401 -28
rect 600 29 606 35
rect 601 6 606 11
rect 483 -40 488 -35
rect 570 -26 575 -21
rect 197 -80 202 -75
rect 197 -89 202 -84
rect 321 -93 326 -88
rect 343 -80 348 -75
rect 347 -92 352 -87
rect 183 -131 188 -126
rect 176 -163 181 -158
rect 169 -172 174 -167
rect 155 -206 160 -201
rect 155 -265 160 -260
rect 169 -256 174 -251
rect 169 -297 174 -292
rect 162 -329 167 -324
rect 155 -338 160 -333
rect 148 -363 153 -358
rect 141 -372 146 -367
rect 141 -438 146 -433
rect 141 -487 146 -482
rect 141 -528 146 -522
rect 155 -430 160 -425
rect 155 -479 160 -474
rect 169 -422 174 -417
rect 197 -131 202 -126
rect 197 -140 202 -135
rect 197 -149 202 -144
rect 197 -163 202 -158
rect 321 -152 326 -147
rect 197 -172 202 -167
rect 197 -181 202 -176
rect 321 -185 326 -180
rect 347 -106 352 -101
rect 396 -99 401 -94
rect 483 -83 488 -78
rect 553 -39 558 -34
rect 594 -41 599 -36
rect 570 -89 575 -84
rect 594 -58 599 -53
rect 483 -131 488 -126
rect 570 -116 575 -111
rect 342 -176 347 -171
rect 342 -185 347 -180
rect 197 -197 202 -192
rect 197 -206 202 -201
rect 321 -210 326 -205
rect 183 -248 188 -243
rect 183 -289 188 -284
rect 347 -197 352 -192
rect 346 -221 352 -215
rect 197 -247 202 -242
rect 197 -256 202 -251
rect 197 -265 202 -260
rect 197 -274 202 -269
rect 321 -277 326 -272
rect 339 -277 344 -272
rect 197 -287 202 -282
rect 197 -296 202 -291
rect 197 -305 202 -300
rect 197 -314 202 -309
rect 197 -329 202 -324
rect 321 -318 326 -313
rect 395 -204 400 -199
rect 483 -172 488 -167
rect 553 -129 558 -124
rect 610 -58 615 -53
rect 664 -66 669 -61
rect 594 -131 599 -126
rect 570 -179 575 -174
rect 594 -148 599 -143
rect 553 -192 558 -187
rect 483 -223 488 -218
rect 570 -205 575 -200
rect 483 -263 488 -258
rect 553 -218 558 -213
rect 610 -139 615 -134
rect 594 -220 599 -215
rect 570 -268 575 -263
rect 594 -237 599 -232
rect 483 -293 488 -288
rect 342 -326 347 -321
rect 197 -338 202 -333
rect 197 -347 202 -342
rect 321 -351 326 -346
rect 342 -335 347 -330
rect 347 -347 352 -342
rect 197 -363 202 -358
rect 197 -372 202 -367
rect 321 -376 326 -371
rect 346 -386 351 -381
rect 197 -422 202 -417
rect 188 -430 193 -425
rect 197 -438 202 -433
rect 197 -447 202 -442
rect 321 -451 326 -446
rect 339 -451 344 -446
rect 177 -479 182 -474
rect 197 -487 202 -482
rect 197 -496 202 -491
rect 321 -500 326 -495
rect 197 -528 202 -523
rect 197 -537 202 -532
rect 321 -541 326 -536
rect 395 -356 400 -351
rect 462 -500 467 -495
rect 570 -293 575 -288
rect 483 -347 488 -342
rect 553 -306 558 -301
rect 610 -220 615 -215
rect 664 -228 669 -223
rect 594 -308 599 -303
rect 570 -356 575 -351
rect 594 -325 599 -320
rect 483 -405 488 -400
rect 570 -382 575 -377
rect 483 -435 488 -430
rect 553 -395 558 -390
rect 610 -301 615 -296
rect 594 -397 599 -392
rect 570 -445 575 -440
rect 594 -414 599 -409
rect 610 -382 615 -377
rect 664 -390 669 -385
rect 610 -463 615 -458
rect 337 -531 342 -526
rect 342 -540 347 -535
rect 339 -549 344 -544
rect 197 -570 202 -564
rect 321 -574 326 -569
rect 347 -561 352 -556
rect 321 -599 326 -594
<< pm12contact >>
rect 162 -197 167 -192
rect 155 -305 160 -300
<< metal2 >>
rect 65 131 176 134
rect 195 131 242 134
rect 78 114 219 117
rect 78 88 183 91
rect -33 74 7 78
rect 78 66 82 88
rect 188 88 235 91
rect 99 75 122 79
rect 118 64 122 75
rect 232 49 235 88
rect 239 56 242 131
rect 239 53 482 56
rect 232 46 470 49
rect 118 15 122 42
rect 220 19 223 44
rect 220 16 347 19
rect 99 11 122 15
rect -34 -6 0 -2
rect 65 -1 162 2
rect 188 -12 197 -8
rect 78 -18 160 -15
rect 326 -16 343 -12
rect 157 -21 160 -18
rect 157 -24 347 -21
rect 401 -32 463 -29
rect 170 -38 392 -35
rect 170 -40 174 -38
rect 78 -44 169 -41
rect 78 -66 82 -44
rect 389 -41 392 -38
rect 389 -44 456 -41
rect 99 -57 122 -53
rect 188 -55 197 -51
rect 118 -68 122 -57
rect 174 -63 197 -59
rect 326 -67 340 -63
rect 336 -75 340 -67
rect 181 -80 197 -76
rect 336 -79 343 -75
rect -33 -87 7 -83
rect 174 -88 197 -84
rect 348 -87 352 -85
rect 118 -117 122 -90
rect 326 -92 347 -88
rect 401 -98 449 -95
rect 133 -105 347 -102
rect 99 -121 122 -117
rect 157 -114 368 -111
rect 65 -136 148 -133
rect 157 -144 160 -114
rect 188 -131 197 -127
rect 174 -139 197 -135
rect 364 -142 367 -114
rect 156 -147 197 -144
rect 78 -153 128 -150
rect -34 -168 -1 -164
rect 156 -175 160 -147
rect 364 -145 442 -142
rect 326 -151 338 -147
rect 181 -163 197 -160
rect 174 -172 197 -168
rect 335 -172 338 -151
rect 78 -179 155 -176
rect 78 -201 82 -179
rect 335 -176 342 -172
rect 347 -176 348 -172
rect 160 -180 197 -176
rect 326 -184 342 -180
rect 347 -184 348 -180
rect 99 -192 122 -188
rect -4 -206 7 -202
rect -4 -245 0 -206
rect 118 -203 122 -192
rect 167 -197 197 -193
rect 160 -205 197 -201
rect 347 -205 351 -197
rect 326 -209 351 -205
rect 396 -207 435 -204
rect -33 -249 0 -245
rect 138 -220 346 -217
rect 118 -252 122 -225
rect 146 -231 366 -228
rect 188 -247 197 -244
rect 99 -256 122 -252
rect 174 -256 197 -252
rect 160 -264 197 -260
rect 65 -268 139 -265
rect 139 -273 197 -269
rect 326 -276 339 -272
rect 78 -285 126 -282
rect 188 -287 197 -284
rect 363 -283 366 -231
rect 432 -276 435 -207
rect 439 -259 442 -145
rect 446 -218 449 -98
rect 453 -167 456 -44
rect 460 -126 463 -32
rect 467 -78 470 46
rect 479 -35 482 53
rect 602 11 605 29
rect 553 -5 610 -2
rect 553 -34 558 -5
rect 575 -25 598 -21
rect 479 -40 483 -35
rect 594 -36 598 -25
rect 607 -57 610 -5
rect 467 -83 483 -78
rect 594 -85 598 -58
rect 669 -66 700 -62
rect 575 -89 598 -85
rect 553 -102 610 -99
rect 553 -124 558 -102
rect 575 -115 598 -111
rect 460 -131 483 -126
rect 594 -126 598 -115
rect 607 -138 610 -102
rect 453 -172 483 -167
rect 594 -175 598 -148
rect 575 -179 598 -175
rect 558 -191 610 -188
rect 481 -200 485 -196
rect 553 -213 558 -192
rect 575 -204 598 -200
rect 594 -215 598 -204
rect 446 -223 483 -218
rect 607 -219 610 -191
rect 669 -228 700 -224
rect 439 -262 483 -259
rect 594 -264 598 -237
rect 575 -268 598 -264
rect 432 -279 482 -276
rect 363 -286 468 -283
rect 174 -296 197 -293
rect 160 -305 197 -301
rect 78 -311 141 -308
rect -34 -329 -1 -325
rect 78 -333 82 -311
rect 146 -312 197 -309
rect 326 -317 338 -313
rect 99 -324 122 -320
rect 335 -322 338 -317
rect 118 -335 122 -324
rect 167 -329 197 -326
rect 335 -326 342 -322
rect 160 -338 197 -334
rect 339 -335 342 -330
rect -4 -346 7 -342
rect -4 -406 0 -346
rect 146 -346 197 -342
rect 339 -346 343 -335
rect 326 -350 343 -346
rect 347 -342 351 -341
rect 465 -343 468 -286
rect 479 -288 482 -279
rect 553 -279 610 -276
rect 479 -292 483 -288
rect 553 -301 558 -279
rect 575 -292 598 -288
rect 594 -303 598 -292
rect 607 -300 610 -279
rect 465 -346 483 -343
rect 118 -384 122 -357
rect 153 -363 197 -359
rect 146 -371 197 -367
rect 347 -371 351 -347
rect 400 -355 466 -352
rect 326 -375 351 -371
rect 99 -387 122 -384
rect 127 -385 346 -382
rect 65 -402 118 -399
rect -33 -410 0 -406
rect 127 -416 130 -385
rect 78 -419 130 -416
rect 138 -397 364 -394
rect 138 -423 141 -397
rect 174 -421 197 -418
rect 128 -426 141 -423
rect 128 -441 131 -426
rect 160 -430 188 -426
rect 361 -431 364 -397
rect 463 -401 466 -355
rect 594 -352 598 -325
rect 575 -356 598 -352
rect 553 -368 610 -365
rect 553 -390 558 -368
rect 575 -381 598 -377
rect 607 -381 610 -368
rect 594 -392 598 -381
rect 669 -390 700 -386
rect 463 -404 483 -401
rect 146 -438 197 -434
rect 361 -434 483 -431
rect 78 -445 127 -442
rect 78 -467 82 -445
rect 132 -446 197 -442
rect 594 -441 598 -414
rect 575 -445 598 -441
rect 326 -450 339 -446
rect 99 -458 122 -454
rect 118 -469 122 -458
rect 615 -462 616 -459
rect 610 -470 615 -463
rect 480 -473 615 -470
rect -3 -478 7 -474
rect 160 -479 177 -475
rect -35 -491 -1 -487
rect 146 -487 197 -483
rect -3 -505 3 -504
rect -7 -508 3 -505
rect -1 -568 3 -508
rect 118 -518 122 -491
rect 132 -495 197 -491
rect 326 -499 339 -495
rect 99 -522 122 -518
rect 146 -528 197 -524
rect 335 -526 339 -499
rect 480 -496 483 -473
rect 610 -496 615 -473
rect 467 -499 483 -496
rect 335 -531 337 -526
rect 132 -536 197 -532
rect 326 -540 342 -536
rect -33 -572 3 -568
rect 132 -569 197 -565
rect 335 -569 339 -544
rect 326 -573 339 -569
rect 347 -594 351 -561
rect 326 -598 351 -594
<< labels >>
rlabel metal1 191 -406 194 130 1 c0
rlabel m2contact 183 87 188 92 1 P0
rlabel m2contact 176 130 181 135 1 G0
rlabel m2contact 162 -2 167 3 1 G1
rlabel m2contact 169 -45 174 -40 1 P1
rlabel m2contact 148 -136 153 -131 1 G2
rlabel m2contact 155 -180 160 -175 1 P2
rlabel m2contact 134 -273 139 -268 1 G3
rlabel m2contact 141 -312 146 -307 1 P3
rlabel m2contact 127 -446 132 -441 1 P4
rlabel metal1 395 -356 399 -302 1 C4
rlabel metal1 396 -99 400 -63 1 C2
rlabel metal1 395 -203 399 -168 1 C3
rlabel polycontact 8 31 12 35 1 a0
rlabel polycontact 8 39 12 43 1 b0
rlabel polycontact 8 -93 12 -89 1 b1
rlabel polycontact 8 -236 12 -232 1 a2
rlabel polycontact 8 -228 12 -224 1 b2
rlabel polycontact 8 -360 12 -356 1 b3
rlabel polycontact 8 -368 12 -364 1 a3
rlabel polycontact 8 -494 12 -490 1 b4
rlabel polycontact 8 -502 12 -498 1 a4
rlabel m2contact 73 -420 78 -415 1 G4_bar
rlabel m2contact 59 -403 65 -398 1 G4
rlabel m2contact 73 -286 78 -281 1 G3_bar
rlabel m2contact 128 -154 133 -149 1 G2_bar
rlabel m2contact 73 -19 78 -14 1 G1_bar
rlabel m2contact 73 113 78 118 1 G0_bar
rlabel metal1 15 -535 19 138 1 vdd
rlabel psubstratepcontact 111 43 115 47 1 gnd
rlabel polycontact 8 -101 12 -97 1 a1
rlabel metal1 111 -613 476 -609 1 gnd
rlabel metal1 209 -604 213 150 1 vdd
rlabel metal1 472 -613 476 -512 7 gnd
rlabel metal1 330 -613 334 0 1 gnd
rlabel ndcontact 257 -16 261 -12 1 t1
rlabel ndcontact 257 -67 261 -63 1 t2
rlabel ndcontact 257 -92 261 -88 1 t3
rlabel ndcontact 256 -151 260 -147 1 t4
rlabel ndcontact 256 -184 260 -180 1 t5
rlabel ndcontact 256 -209 260 -205 1 t6
rlabel ndcontact 256 -276 260 -272 1 t7
rlabel ndcontact 256 -317 260 -313 1 t8
rlabel ndcontact 256 -350 260 -346 1 t9
rlabel ndcontact 256 -375 260 -371 1 t10
rlabel ndcontact 256 -450 260 -446 1 t11
rlabel ndcontact 256 -499 260 -495 1 t12
rlabel ndcontact 256 -540 260 -536 1 t13
rlabel ndcontact 256 -573 260 -569 1 t14
rlabel ndcontact 256 -598 260 -594 1 t15
rlabel metal1 -15 -2 -11 1 7 gnd
rlabel m2contact -37 74 -33 77 5 Q
rlabel polycontact -39 63 -35 67 7 Q_bar
rlabel polycontact -38 39 -34 43 7 Y
rlabel polycontact -44 18 -40 22 7 X
rlabel pdiffusion -68 6 -48 10 7 l1
rlabel ndiffusion -30 22 -20 26 7 l2
rlabel ndiffusion -30 46 -20 50 7 l3
rlabel ndiffusion -30 127 -20 131 7 l3
rlabel ndiffusion -30 103 -20 107 7 l2
rlabel pdiffusion -68 87 -48 91 7 l1
rlabel polycontact -44 99 -40 103 7 X
rlabel polycontact -38 120 -34 124 7 Y
rlabel polycontact -39 144 -35 148 7 Q_bar
rlabel metal1 -37 155 -33 165 5 Q
rlabel metal1 -15 83 -11 161 7 gnd
rlabel metal1 -80 -8 -76 80 7 vdd
rlabel metal1 -80 73 -76 161 7 vdd
rlabel polycontact -87 10 -83 14 3 clk
rlabel polycontact -87 2 -83 6 3 D
rlabel polycontact -87 83 -83 87 3 D
rlabel polycontact -87 91 -83 95 3 clk
rlabel metal1 -15 -163 -11 -77 7 gnd
rlabel m2contact -37 -87 -33 -84 5 Q
rlabel polycontact -39 -98 -35 -94 7 Q_bar
rlabel polycontact -38 -122 -34 -118 7 Y
rlabel polycontact -44 -143 -40 -139 7 X
rlabel ndiffusion -30 -139 -20 -135 7 l2
rlabel ndiffusion -30 -115 -20 -111 7 l3
rlabel ndiffusion -30 -34 -20 -30 7 l3
rlabel ndiffusion -30 -58 -20 -54 7 l2
rlabel pdiffusion -68 -74 -48 -70 7 l1
rlabel polycontact -44 -62 -40 -58 7 X
rlabel polycontact -38 -41 -34 -37 7 Y
rlabel polycontact -39 -17 -35 -13 7 Q_bar
rlabel metal1 -15 -78 -11 1 7 gnd
rlabel metal1 -80 -169 -76 -81 7 vdd
rlabel metal1 -80 -88 -76 0 7 vdd
rlabel polycontact -87 -78 -83 -74 3 D
rlabel polycontact -87 -70 -83 -66 3 clk
rlabel polycontact -87 -159 -83 -155 3 D
rlabel polycontact -87 -151 -83 -147 3 clk
rlabel pdiffusion -68 -155 -48 -151 7 l1
rlabel metal1 -15 -325 -11 -239 7 gnd
rlabel m2contact -37 -249 -33 -246 5 Q
rlabel polycontact -39 -260 -35 -256 7 Q_bar
rlabel polycontact -38 -284 -34 -280 7 Y
rlabel polycontact -44 -305 -40 -301 7 X
rlabel pdiffusion -68 -317 -48 -313 7 l1
rlabel ndiffusion -30 -301 -20 -297 7 l2
rlabel ndiffusion -30 -277 -20 -273 7 l3
rlabel ndiffusion -30 -196 -20 -192 7 l3
rlabel ndiffusion -30 -220 -20 -216 7 l2
rlabel pdiffusion -68 -236 -48 -232 7 l1
rlabel polycontact -44 -224 -40 -220 7 X
rlabel polycontact -38 -203 -34 -199 7 Y
rlabel polycontact -39 -179 -35 -175 7 Q_bar
rlabel metal1 -15 -240 -11 -161 7 gnd
rlabel metal1 -80 -331 -76 -243 7 vdd
rlabel metal1 -80 -250 -76 -162 7 vdd
rlabel polycontact -87 -313 -83 -309 3 clk
rlabel polycontact -87 -321 -83 -317 3 D
rlabel polycontact -87 -240 -83 -236 3 D
rlabel polycontact -87 -232 -83 -228 3 clk
rlabel polycontact -87 -393 -83 -389 3 clk
rlabel polycontact -87 -401 -83 -397 3 D
rlabel polycontact -87 -482 -83 -478 3 D
rlabel metal1 -80 -411 -76 -323 7 vdd
rlabel metal1 -80 -492 -76 -404 7 vdd
rlabel metal1 -15 -401 -11 -322 7 gnd
rlabel polycontact -39 -340 -35 -336 7 Q_bar
rlabel polycontact -38 -364 -34 -360 7 Y
rlabel polycontact -44 -385 -40 -381 7 X
rlabel pdiffusion -68 -397 -48 -393 7 l1
rlabel ndiffusion -30 -381 -20 -377 7 l2
rlabel ndiffusion -30 -357 -20 -353 7 l3
rlabel ndiffusion -30 -438 -20 -434 7 l3
rlabel ndiffusion -30 -462 -20 -458 7 l2
rlabel pdiffusion -68 -478 -48 -474 7 l1
rlabel polycontact -44 -466 -40 -462 7 X
rlabel polycontact -38 -445 -34 -441 7 Y
rlabel polycontact -39 -421 -35 -417 7 Q_bar
rlabel m2contact -37 -410 -33 -407 5 Q
rlabel metal1 -15 -486 -11 -400 7 gnd
rlabel metal1 -15 -648 -11 -562 7 gnd
rlabel m2contact -37 -572 -33 -569 5 Q
rlabel polycontact -39 -583 -35 -579 7 Q_bar
rlabel polycontact -38 -607 -34 -603 7 Y
rlabel polycontact -44 -628 -40 -624 7 X
rlabel pdiffusion -68 -640 -48 -636 7 l1
rlabel ndiffusion -30 -624 -20 -620 7 l2
rlabel ndiffusion -30 -600 -20 -596 7 l3
rlabel ndiffusion -30 -519 -20 -515 7 l3
rlabel ndiffusion -30 -543 -20 -539 7 l2
rlabel pdiffusion -68 -559 -48 -555 7 l1
rlabel polycontact -44 -547 -40 -543 7 X
rlabel polycontact -38 -526 -34 -522 7 Y
rlabel polycontact -39 -502 -35 -498 7 Q_bar
rlabel metal1 -15 -563 -11 -484 7 gnd
rlabel metal1 -80 -654 -76 -566 7 vdd
rlabel metal1 -80 -573 -76 -485 7 vdd
rlabel polycontact -87 -636 -83 -632 3 clk
rlabel polycontact -87 -644 -83 -640 3 D
rlabel polycontact -87 -563 -83 -559 3 D
rlabel polycontact -87 -555 -83 -551 3 clk
rlabel metal1 397 -34 401 -33 1 C1
rlabel metal1 491 -459 495 -363 7 vdd
rlabel metal1 587 -459 591 -363 7 gnd
rlabel metal1 498 -429 501 -393 7 l4
rlabel polycontact 484 -417 488 -413 3 B
rlabel polycontact 484 -425 488 -421 7 A
rlabel polycontact 594 -409 598 -405 7 A_bar
rlabel polycontact 594 -401 598 -397 7 B_bar
rlabel ndiffusion 561 -421 581 -417 7 l1
rlabel ndiffusion 561 -405 581 -401 7 l2
rlabel pdiffusion 505 -413 545 -409 7 l3
rlabel metal1 491 -370 495 -274 7 vdd
rlabel metal1 587 -370 591 -274 7 gnd
rlabel metal1 498 -340 501 -304 7 l4
rlabel polycontact 484 -328 488 -324 3 B
rlabel polycontact 484 -336 488 -332 7 A
rlabel polycontact 594 -320 598 -316 7 A_bar
rlabel polycontact 594 -312 598 -308 7 B_bar
rlabel ndiffusion 561 -332 581 -328 7 l1
rlabel ndiffusion 561 -316 581 -312 7 l2
rlabel pdiffusion 505 -324 545 -320 7 l3
rlabel metal1 491 -282 495 -186 7 vdd
rlabel metal1 587 -282 591 -186 7 gnd
rlabel metal1 498 -252 501 -216 7 l4
rlabel polycontact 484 -240 488 -236 3 B
rlabel polycontact 484 -248 488 -244 7 A
rlabel polycontact 594 -232 598 -228 7 A_bar
rlabel polycontact 594 -224 598 -220 7 B_bar
rlabel ndiffusion 561 -244 581 -240 7 l1
rlabel ndiffusion 561 -228 581 -224 7 l2
rlabel pdiffusion 505 -236 545 -232 7 l3
rlabel metal1 498 -163 501 -127 7 l4
rlabel metal1 491 -193 495 -97 7 vdd
rlabel polycontact 484 -151 488 -147 3 B
rlabel polycontact 484 -159 488 -155 7 A
rlabel polycontact 594 -143 598 -139 7 A_bar
rlabel metal1 587 -193 591 -97 7 gnd
rlabel polycontact 594 -135 598 -131 7 B_bar
rlabel ndiffusion 561 -155 581 -151 7 l1
rlabel ndiffusion 561 -139 581 -135 7 l2
rlabel pdiffusion 505 -147 545 -143 7 l3
rlabel pdiffusion 505 -57 545 -53 7 l3
rlabel ndiffusion 561 -49 581 -45 7 l2
rlabel ndiffusion 561 -65 581 -61 7 l1
rlabel polycontact 594 -45 598 -41 7 B_bar
rlabel polycontact 594 -53 598 -49 7 A_bar
rlabel polycontact 484 -69 488 -65 7 A
rlabel polycontact 484 -61 488 -57 3 B
rlabel metal1 498 -73 501 -37 7 l4
rlabel metal1 587 -103 591 -7 7 gnd
rlabel metal1 491 -103 495 -7 7 vdd
rlabel polycontact 615 -373 619 -369 3 clk
rlabel polycontact 615 -381 619 -377 3 D
rlabel polycontact 615 -462 619 -458 3 D
rlabel polycontact 615 -454 619 -450 3 clk
rlabel metal1 622 -391 626 -303 7 vdd
rlabel metal1 622 -472 626 -384 7 vdd
rlabel metal1 687 -381 691 -302 7 gnd
rlabel polycontact 663 -320 667 -316 7 Q_bar
rlabel polycontact 664 -344 668 -340 7 Y
rlabel polycontact 658 -365 662 -361 7 X
rlabel pdiffusion 634 -377 654 -373 7 l1
rlabel ndiffusion 672 -361 682 -357 7 l2
rlabel ndiffusion 672 -337 682 -333 7 l3
rlabel ndiffusion 672 -418 682 -414 7 l3
rlabel ndiffusion 672 -442 682 -438 7 l2
rlabel pdiffusion 634 -458 654 -454 7 l1
rlabel polycontact 658 -446 662 -442 7 X
rlabel polycontact 664 -425 668 -421 7 Y
rlabel polycontact 663 -401 667 -397 7 Q_bar
rlabel m2contact 665 -390 669 -387 5 Q
rlabel metal1 687 -466 691 -380 7 gnd
rlabel metal1 622 -310 626 -222 7 vdd
rlabel metal1 687 -304 691 -218 7 gnd
rlabel m2contact 665 -228 669 -225 5 Q
rlabel polycontact 663 -239 667 -235 7 Q_bar
rlabel polycontact 664 -263 668 -259 7 Y
rlabel polycontact 658 -284 662 -280 7 X
rlabel pdiffusion 634 -296 654 -292 7 l1
rlabel ndiffusion 672 -280 682 -276 7 l2
rlabel ndiffusion 672 -256 682 -252 7 l3
rlabel ndiffusion 672 -175 682 -171 7 l3
rlabel ndiffusion 672 -199 682 -195 7 l2
rlabel pdiffusion 634 -215 654 -211 7 l1
rlabel polycontact 658 -203 662 -199 7 X
rlabel polycontact 664 -182 668 -178 7 Y
rlabel polycontact 663 -158 667 -154 7 Q_bar
rlabel metal1 687 -219 691 -140 7 gnd
rlabel metal1 622 -229 626 -141 7 vdd
rlabel polycontact 615 -292 619 -288 3 clk
rlabel polycontact 615 -219 619 -215 3 D
rlabel polycontact 615 -211 619 -207 3 clk
rlabel metal1 622 -148 626 -60 7 vdd
rlabel polycontact 615 -49 619 -45 3 clk
rlabel polycontact 615 -57 619 -53 3 D
rlabel polycontact 615 -138 619 -134 3 D
rlabel polycontact 615 -130 619 -126 3 clk
rlabel metal1 622 -67 626 21 7 vdd
rlabel metal1 687 -57 691 19 7 gnd
rlabel polycontact 663 4 667 8 7 Q_bar
rlabel polycontact 664 -20 668 -16 7 Y
rlabel polycontact 658 -41 662 -37 7 X
rlabel pdiffusion 634 -53 654 -49 7 l1
rlabel ndiffusion 672 -37 682 -33 7 l2
rlabel ndiffusion 672 -13 682 -9 7 l3
rlabel ndiffusion 672 -94 682 -90 7 l3
rlabel ndiffusion 672 -118 682 -114 7 l2
rlabel pdiffusion 634 -134 654 -130 7 l1
rlabel polycontact 658 -122 662 -118 7 X
rlabel polycontact 664 -101 668 -97 7 Y
rlabel polycontact 663 -77 667 -73 7 Q_bar
rlabel m2contact 665 -66 669 -63 5 Q
rlabel metal1 687 -142 691 -56 7 gnd
rlabel metal1 276 104 362 108 1 gnd
rlabel metal1 276 126 286 130 3 Q
rlabel polycontact 293 128 297 132 1 Q_bar
rlabel polycontact 317 127 321 131 1 Y
rlabel polycontact 338 133 342 137 1 X
rlabel pdiffusion 350 141 354 161 1 l1
rlabel ndiffusion 334 113 338 123 1 l2
rlabel ndiffusion 310 113 314 123 1 l3
rlabel polycontact 346 176 350 180 5 clk
rlabel polycontact 354 176 358 180 5 D
<< end >>
