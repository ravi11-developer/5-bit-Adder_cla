magic
tech scmos
timestamp 1764674403
<< nwell >>
rect -448 723 -422 757
rect -609 668 -485 705
rect -392 655 -330 698
rect -611 566 -487 603
rect -315 559 -255 617
rect -449 511 -423 545
rect -448 223 -422 257
rect -609 168 -485 205
rect -392 155 -330 198
rect -611 66 -487 103
rect -315 59 -255 117
rect -449 11 -423 45
rect -449 -224 -423 -190
rect -611 -279 -487 -242
rect -393 -292 -331 -249
rect -612 -381 -488 -344
rect -316 -388 -256 -330
rect -450 -436 -424 -402
rect -447 -685 -421 -651
rect -613 -740 -489 -703
rect -391 -753 -329 -710
rect -611 -843 -487 -806
rect -314 -849 -254 -791
rect -448 -897 -422 -863
rect -446 -1039 -420 -1005
rect -611 -1090 -487 -1053
rect -390 -1107 -328 -1064
rect -610 -1200 -486 -1163
rect -313 -1203 -253 -1145
rect -88 -1211 -24 -1186
rect -447 -1251 -421 -1217
rect -88 -1244 -25 -1211
rect -88 -1245 -51 -1244
<< ntransistor >>
rect -436 700 -434 710
rect -598 643 -596 653
rect -563 643 -561 653
rect -551 643 -549 653
rect -530 643 -528 653
rect -518 643 -516 653
rect -498 643 -496 653
rect -381 616 -379 636
rect -369 616 -367 636
rect -344 632 -342 642
rect -600 541 -598 551
rect -565 541 -563 551
rect -553 541 -551 551
rect -532 541 -530 551
rect -520 541 -518 551
rect -500 541 -498 551
rect -304 500 -302 520
rect -292 500 -290 520
rect -280 500 -278 520
rect -268 500 -266 520
rect -437 488 -435 498
rect -436 200 -434 210
rect -598 143 -596 153
rect -563 143 -561 153
rect -551 143 -549 153
rect -530 143 -528 153
rect -518 143 -516 153
rect -498 143 -496 153
rect -381 116 -379 136
rect -369 116 -367 136
rect -344 132 -342 142
rect -600 41 -598 51
rect -565 41 -563 51
rect -553 41 -551 51
rect -532 41 -530 51
rect -520 41 -518 51
rect -500 41 -498 51
rect -304 0 -302 20
rect -292 0 -290 20
rect -280 0 -278 20
rect -268 0 -266 20
rect -437 -12 -435 -2
rect -437 -247 -435 -237
rect -600 -304 -598 -294
rect -565 -304 -563 -294
rect -553 -304 -551 -294
rect -532 -304 -530 -294
rect -520 -304 -518 -294
rect -500 -304 -498 -294
rect -382 -331 -380 -311
rect -370 -331 -368 -311
rect -345 -315 -343 -305
rect -601 -406 -599 -396
rect -566 -406 -564 -396
rect -554 -406 -552 -396
rect -533 -406 -531 -396
rect -521 -406 -519 -396
rect -501 -406 -499 -396
rect -305 -447 -303 -427
rect -293 -447 -291 -427
rect -281 -447 -279 -427
rect -269 -447 -267 -427
rect -438 -459 -436 -449
rect -435 -708 -433 -698
rect -602 -765 -600 -755
rect -567 -765 -565 -755
rect -555 -765 -553 -755
rect -534 -765 -532 -755
rect -522 -765 -520 -755
rect -502 -765 -500 -755
rect -380 -792 -378 -772
rect -368 -792 -366 -772
rect -343 -776 -341 -766
rect -600 -868 -598 -858
rect -565 -868 -563 -858
rect -553 -868 -551 -858
rect -532 -868 -530 -858
rect -520 -868 -518 -858
rect -500 -868 -498 -858
rect -303 -908 -301 -888
rect -291 -908 -289 -888
rect -279 -908 -277 -888
rect -267 -908 -265 -888
rect -436 -920 -434 -910
rect -434 -1062 -432 -1052
rect -600 -1115 -598 -1105
rect -565 -1115 -563 -1105
rect -553 -1115 -551 -1105
rect -532 -1115 -530 -1105
rect -520 -1115 -518 -1105
rect -500 -1115 -498 -1105
rect -379 -1146 -377 -1126
rect -367 -1146 -365 -1126
rect -342 -1130 -340 -1120
rect -599 -1225 -597 -1215
rect -564 -1225 -562 -1215
rect -552 -1225 -550 -1215
rect -531 -1225 -529 -1215
rect -519 -1225 -517 -1215
rect -499 -1225 -497 -1215
rect -302 -1262 -300 -1242
rect -290 -1262 -288 -1242
rect -278 -1262 -276 -1242
rect -266 -1262 -264 -1242
rect -435 -1274 -433 -1264
rect -76 -1273 -74 -1263
rect -64 -1273 -62 -1263
rect -39 -1267 -37 -1257
<< ptransistor >>
rect -436 730 -434 750
rect -598 674 -596 694
rect -586 674 -584 694
rect -563 674 -561 694
rect -530 674 -528 694
rect -498 674 -496 694
rect -381 661 -379 681
rect -369 661 -367 681
rect -344 662 -342 682
rect -600 572 -598 592
rect -588 572 -586 592
rect -565 572 -563 592
rect -532 572 -530 592
rect -500 572 -498 592
rect -304 565 -302 605
rect -292 565 -290 605
rect -280 565 -278 605
rect -268 565 -266 605
rect -437 518 -435 538
rect -436 230 -434 250
rect -598 174 -596 194
rect -586 174 -584 194
rect -563 174 -561 194
rect -530 174 -528 194
rect -498 174 -496 194
rect -381 161 -379 181
rect -369 161 -367 181
rect -344 162 -342 182
rect -600 72 -598 92
rect -588 72 -586 92
rect -565 72 -563 92
rect -532 72 -530 92
rect -500 72 -498 92
rect -304 65 -302 105
rect -292 65 -290 105
rect -280 65 -278 105
rect -268 65 -266 105
rect -437 18 -435 38
rect -437 -217 -435 -197
rect -600 -273 -598 -253
rect -588 -273 -586 -253
rect -565 -273 -563 -253
rect -532 -273 -530 -253
rect -500 -273 -498 -253
rect -382 -286 -380 -266
rect -370 -286 -368 -266
rect -345 -285 -343 -265
rect -601 -375 -599 -355
rect -589 -375 -587 -355
rect -566 -375 -564 -355
rect -533 -375 -531 -355
rect -501 -375 -499 -355
rect -305 -382 -303 -342
rect -293 -382 -291 -342
rect -281 -382 -279 -342
rect -269 -382 -267 -342
rect -438 -429 -436 -409
rect -435 -678 -433 -658
rect -602 -734 -600 -714
rect -590 -734 -588 -714
rect -567 -734 -565 -714
rect -534 -734 -532 -714
rect -502 -734 -500 -714
rect -380 -747 -378 -727
rect -368 -747 -366 -727
rect -343 -746 -341 -726
rect -600 -837 -598 -817
rect -588 -837 -586 -817
rect -565 -837 -563 -817
rect -532 -837 -530 -817
rect -500 -837 -498 -817
rect -303 -843 -301 -803
rect -291 -843 -289 -803
rect -279 -843 -277 -803
rect -267 -843 -265 -803
rect -436 -890 -434 -870
rect -434 -1032 -432 -1012
rect -600 -1084 -598 -1064
rect -588 -1084 -586 -1064
rect -565 -1084 -563 -1064
rect -532 -1084 -530 -1064
rect -500 -1084 -498 -1064
rect -379 -1101 -377 -1081
rect -367 -1101 -365 -1081
rect -342 -1100 -340 -1080
rect -599 -1194 -597 -1174
rect -587 -1194 -585 -1174
rect -564 -1194 -562 -1174
rect -531 -1194 -529 -1174
rect -499 -1194 -497 -1174
rect -302 -1197 -300 -1157
rect -290 -1197 -288 -1157
rect -278 -1197 -276 -1157
rect -266 -1197 -264 -1157
rect -435 -1244 -433 -1224
rect -76 -1239 -74 -1199
rect -64 -1239 -62 -1199
rect -39 -1237 -37 -1217
<< ndiffusion >>
rect -437 700 -436 710
rect -434 700 -433 710
rect -599 643 -598 653
rect -596 643 -595 653
rect -564 643 -563 653
rect -561 643 -551 653
rect -549 643 -548 653
rect -531 643 -530 653
rect -528 643 -518 653
rect -516 643 -515 653
rect -499 643 -498 653
rect -496 643 -495 653
rect -382 616 -381 636
rect -379 616 -369 636
rect -367 616 -366 636
rect -345 632 -344 642
rect -342 632 -341 642
rect -601 541 -600 551
rect -598 541 -597 551
rect -566 541 -565 551
rect -563 541 -553 551
rect -551 541 -550 551
rect -533 541 -532 551
rect -530 541 -520 551
rect -518 541 -517 551
rect -501 541 -500 551
rect -498 541 -497 551
rect -305 500 -304 520
rect -302 500 -292 520
rect -290 500 -289 520
rect -281 500 -280 520
rect -278 500 -268 520
rect -266 500 -265 520
rect -438 488 -437 498
rect -435 488 -434 498
rect -437 200 -436 210
rect -434 200 -433 210
rect -599 143 -598 153
rect -596 143 -595 153
rect -564 143 -563 153
rect -561 143 -551 153
rect -549 143 -548 153
rect -531 143 -530 153
rect -528 143 -518 153
rect -516 143 -515 153
rect -499 143 -498 153
rect -496 143 -495 153
rect -382 116 -381 136
rect -379 116 -369 136
rect -367 116 -366 136
rect -345 132 -344 142
rect -342 132 -341 142
rect -601 41 -600 51
rect -598 41 -597 51
rect -566 41 -565 51
rect -563 41 -553 51
rect -551 41 -550 51
rect -533 41 -532 51
rect -530 41 -520 51
rect -518 41 -517 51
rect -501 41 -500 51
rect -498 41 -497 51
rect -305 0 -304 20
rect -302 0 -292 20
rect -290 0 -289 20
rect -281 0 -280 20
rect -278 0 -268 20
rect -266 0 -265 20
rect -438 -12 -437 -2
rect -435 -12 -434 -2
rect -438 -247 -437 -237
rect -435 -247 -434 -237
rect -601 -304 -600 -294
rect -598 -304 -597 -294
rect -566 -304 -565 -294
rect -563 -304 -553 -294
rect -551 -304 -550 -294
rect -533 -304 -532 -294
rect -530 -304 -520 -294
rect -518 -304 -517 -294
rect -501 -304 -500 -294
rect -498 -304 -497 -294
rect -383 -331 -382 -311
rect -380 -331 -370 -311
rect -368 -331 -367 -311
rect -346 -315 -345 -305
rect -343 -315 -342 -305
rect -602 -406 -601 -396
rect -599 -406 -598 -396
rect -567 -406 -566 -396
rect -564 -406 -554 -396
rect -552 -406 -551 -396
rect -534 -406 -533 -396
rect -531 -406 -521 -396
rect -519 -406 -518 -396
rect -502 -406 -501 -396
rect -499 -406 -498 -396
rect -306 -447 -305 -427
rect -303 -447 -293 -427
rect -291 -447 -290 -427
rect -282 -447 -281 -427
rect -279 -447 -269 -427
rect -267 -447 -266 -427
rect -439 -459 -438 -449
rect -436 -459 -435 -449
rect -436 -708 -435 -698
rect -433 -708 -432 -698
rect -603 -765 -602 -755
rect -600 -765 -599 -755
rect -568 -765 -567 -755
rect -565 -765 -555 -755
rect -553 -765 -552 -755
rect -535 -765 -534 -755
rect -532 -765 -522 -755
rect -520 -765 -519 -755
rect -503 -765 -502 -755
rect -500 -765 -499 -755
rect -381 -792 -380 -772
rect -378 -792 -368 -772
rect -366 -792 -365 -772
rect -344 -776 -343 -766
rect -341 -776 -340 -766
rect -601 -868 -600 -858
rect -598 -868 -597 -858
rect -566 -868 -565 -858
rect -563 -868 -553 -858
rect -551 -868 -550 -858
rect -533 -868 -532 -858
rect -530 -868 -520 -858
rect -518 -868 -517 -858
rect -501 -868 -500 -858
rect -498 -868 -497 -858
rect -304 -908 -303 -888
rect -301 -908 -291 -888
rect -289 -908 -288 -888
rect -280 -908 -279 -888
rect -277 -908 -267 -888
rect -265 -908 -264 -888
rect -437 -920 -436 -910
rect -434 -920 -433 -910
rect -435 -1062 -434 -1052
rect -432 -1062 -431 -1052
rect -601 -1115 -600 -1105
rect -598 -1115 -597 -1105
rect -566 -1115 -565 -1105
rect -563 -1115 -553 -1105
rect -551 -1115 -550 -1105
rect -533 -1115 -532 -1105
rect -530 -1115 -520 -1105
rect -518 -1115 -517 -1105
rect -501 -1115 -500 -1105
rect -498 -1115 -497 -1105
rect -380 -1146 -379 -1126
rect -377 -1146 -367 -1126
rect -365 -1146 -364 -1126
rect -343 -1130 -342 -1120
rect -340 -1130 -339 -1120
rect -600 -1225 -599 -1215
rect -597 -1225 -596 -1215
rect -565 -1225 -564 -1215
rect -562 -1225 -552 -1215
rect -550 -1225 -549 -1215
rect -532 -1225 -531 -1215
rect -529 -1225 -519 -1215
rect -517 -1225 -516 -1215
rect -500 -1225 -499 -1215
rect -497 -1225 -496 -1215
rect -303 -1262 -302 -1242
rect -300 -1262 -290 -1242
rect -288 -1262 -287 -1242
rect -279 -1262 -278 -1242
rect -276 -1262 -266 -1242
rect -264 -1262 -263 -1242
rect -436 -1274 -435 -1264
rect -433 -1274 -432 -1264
rect -77 -1273 -76 -1263
rect -74 -1273 -73 -1263
rect -65 -1273 -64 -1263
rect -62 -1273 -61 -1263
rect -40 -1267 -39 -1257
rect -37 -1267 -36 -1257
<< pdiffusion >>
rect -437 730 -436 750
rect -434 730 -433 750
rect -599 674 -598 694
rect -596 674 -586 694
rect -584 674 -583 694
rect -564 674 -563 694
rect -561 674 -560 694
rect -531 674 -530 694
rect -528 674 -527 694
rect -499 674 -498 694
rect -496 674 -495 694
rect -382 661 -381 681
rect -379 661 -378 681
rect -370 661 -369 681
rect -367 661 -366 681
rect -345 662 -344 682
rect -342 662 -341 682
rect -601 572 -600 592
rect -598 572 -588 592
rect -586 572 -585 592
rect -566 572 -565 592
rect -563 572 -562 592
rect -533 572 -532 592
rect -530 572 -529 592
rect -501 572 -500 592
rect -498 572 -497 592
rect -305 565 -304 605
rect -302 565 -292 605
rect -290 565 -289 605
rect -281 565 -280 605
rect -278 565 -268 605
rect -266 565 -265 605
rect -438 518 -437 538
rect -435 518 -434 538
rect -437 230 -436 250
rect -434 230 -433 250
rect -599 174 -598 194
rect -596 174 -586 194
rect -584 174 -583 194
rect -564 174 -563 194
rect -561 174 -560 194
rect -531 174 -530 194
rect -528 174 -527 194
rect -499 174 -498 194
rect -496 174 -495 194
rect -382 161 -381 181
rect -379 161 -378 181
rect -370 161 -369 181
rect -367 161 -366 181
rect -345 162 -344 182
rect -342 162 -341 182
rect -601 72 -600 92
rect -598 72 -588 92
rect -586 72 -585 92
rect -566 72 -565 92
rect -563 72 -562 92
rect -533 72 -532 92
rect -530 72 -529 92
rect -501 72 -500 92
rect -498 72 -497 92
rect -305 65 -304 105
rect -302 65 -292 105
rect -290 65 -289 105
rect -281 65 -280 105
rect -278 65 -268 105
rect -266 65 -265 105
rect -438 18 -437 38
rect -435 18 -434 38
rect -438 -217 -437 -197
rect -435 -217 -434 -197
rect -601 -273 -600 -253
rect -598 -273 -588 -253
rect -586 -273 -585 -253
rect -566 -273 -565 -253
rect -563 -273 -562 -253
rect -533 -273 -532 -253
rect -530 -273 -529 -253
rect -501 -273 -500 -253
rect -498 -273 -497 -253
rect -383 -286 -382 -266
rect -380 -286 -379 -266
rect -371 -286 -370 -266
rect -368 -286 -367 -266
rect -346 -285 -345 -265
rect -343 -285 -342 -265
rect -602 -375 -601 -355
rect -599 -375 -589 -355
rect -587 -375 -586 -355
rect -567 -375 -566 -355
rect -564 -375 -563 -355
rect -534 -375 -533 -355
rect -531 -375 -530 -355
rect -502 -375 -501 -355
rect -499 -375 -498 -355
rect -306 -382 -305 -342
rect -303 -382 -293 -342
rect -291 -382 -290 -342
rect -282 -382 -281 -342
rect -279 -382 -269 -342
rect -267 -382 -266 -342
rect -439 -429 -438 -409
rect -436 -429 -435 -409
rect -436 -678 -435 -658
rect -433 -678 -432 -658
rect -603 -734 -602 -714
rect -600 -734 -590 -714
rect -588 -734 -587 -714
rect -568 -734 -567 -714
rect -565 -734 -564 -714
rect -535 -734 -534 -714
rect -532 -734 -531 -714
rect -503 -734 -502 -714
rect -500 -734 -499 -714
rect -381 -747 -380 -727
rect -378 -747 -377 -727
rect -369 -747 -368 -727
rect -366 -747 -365 -727
rect -344 -746 -343 -726
rect -341 -746 -340 -726
rect -601 -837 -600 -817
rect -598 -837 -588 -817
rect -586 -837 -585 -817
rect -566 -837 -565 -817
rect -563 -837 -562 -817
rect -533 -837 -532 -817
rect -530 -837 -529 -817
rect -501 -837 -500 -817
rect -498 -837 -497 -817
rect -304 -843 -303 -803
rect -301 -843 -291 -803
rect -289 -843 -288 -803
rect -280 -843 -279 -803
rect -277 -843 -267 -803
rect -265 -843 -264 -803
rect -437 -890 -436 -870
rect -434 -890 -433 -870
rect -435 -1032 -434 -1012
rect -432 -1032 -431 -1012
rect -601 -1084 -600 -1064
rect -598 -1084 -588 -1064
rect -586 -1084 -585 -1064
rect -566 -1084 -565 -1064
rect -563 -1084 -562 -1064
rect -533 -1084 -532 -1064
rect -530 -1084 -529 -1064
rect -501 -1084 -500 -1064
rect -498 -1084 -497 -1064
rect -380 -1101 -379 -1081
rect -377 -1101 -376 -1081
rect -368 -1101 -367 -1081
rect -365 -1101 -364 -1081
rect -343 -1100 -342 -1080
rect -340 -1100 -339 -1080
rect -600 -1194 -599 -1174
rect -597 -1194 -587 -1174
rect -585 -1194 -584 -1174
rect -565 -1194 -564 -1174
rect -562 -1194 -561 -1174
rect -532 -1194 -531 -1174
rect -529 -1194 -528 -1174
rect -500 -1194 -499 -1174
rect -497 -1194 -496 -1174
rect -303 -1197 -302 -1157
rect -300 -1197 -290 -1157
rect -288 -1197 -287 -1157
rect -279 -1197 -278 -1157
rect -276 -1197 -266 -1157
rect -264 -1197 -263 -1157
rect -436 -1244 -435 -1224
rect -433 -1244 -432 -1224
rect -77 -1239 -76 -1199
rect -74 -1239 -64 -1199
rect -62 -1239 -61 -1199
rect -40 -1237 -39 -1217
rect -37 -1237 -36 -1217
<< ndcontact >>
rect -441 700 -437 710
rect -433 700 -429 710
rect -603 643 -599 653
rect -595 643 -591 653
rect -568 643 -564 653
rect -548 643 -544 653
rect -535 643 -531 653
rect -515 643 -511 653
rect -503 643 -499 653
rect -495 643 -491 653
rect -386 616 -382 636
rect -366 616 -362 636
rect -349 632 -345 642
rect -341 632 -337 642
rect -386 607 -382 611
rect -376 607 -372 611
rect -366 607 -362 611
rect -344 607 -340 611
rect -605 541 -601 551
rect -597 541 -593 551
rect -570 541 -566 551
rect -550 541 -546 551
rect -537 541 -533 551
rect -517 541 -513 551
rect -505 541 -501 551
rect -497 541 -493 551
rect -309 500 -305 520
rect -289 500 -281 520
rect -265 500 -261 520
rect -442 488 -438 498
rect -434 488 -430 498
rect -441 200 -437 210
rect -433 200 -429 210
rect -603 143 -599 153
rect -595 143 -591 153
rect -568 143 -564 153
rect -548 143 -544 153
rect -535 143 -531 153
rect -515 143 -511 153
rect -503 143 -499 153
rect -495 143 -491 153
rect -386 116 -382 136
rect -366 116 -362 136
rect -349 132 -345 142
rect -341 132 -337 142
rect -386 107 -382 111
rect -376 107 -372 111
rect -366 107 -362 111
rect -344 107 -340 111
rect -605 41 -601 51
rect -597 41 -593 51
rect -570 41 -566 51
rect -550 41 -546 51
rect -537 41 -533 51
rect -517 41 -513 51
rect -505 41 -501 51
rect -497 41 -493 51
rect -309 0 -305 20
rect -289 0 -281 20
rect -265 0 -261 20
rect -442 -12 -438 -2
rect -434 -12 -430 -2
rect -442 -247 -438 -237
rect -434 -247 -430 -237
rect -605 -304 -601 -294
rect -597 -304 -593 -294
rect -570 -304 -566 -294
rect -550 -304 -546 -294
rect -537 -304 -533 -294
rect -517 -304 -513 -294
rect -505 -304 -501 -294
rect -497 -304 -493 -294
rect -387 -331 -383 -311
rect -367 -331 -363 -311
rect -350 -315 -346 -305
rect -342 -315 -338 -305
rect -387 -340 -383 -336
rect -377 -340 -373 -336
rect -367 -340 -363 -336
rect -345 -340 -341 -336
rect -606 -406 -602 -396
rect -598 -406 -594 -396
rect -571 -406 -567 -396
rect -551 -406 -547 -396
rect -538 -406 -534 -396
rect -518 -406 -514 -396
rect -506 -406 -502 -396
rect -498 -406 -494 -396
rect -310 -447 -306 -427
rect -290 -447 -282 -427
rect -266 -447 -262 -427
rect -443 -459 -439 -449
rect -435 -459 -431 -449
rect -440 -708 -436 -698
rect -432 -708 -428 -698
rect -607 -765 -603 -755
rect -599 -765 -595 -755
rect -572 -765 -568 -755
rect -552 -765 -548 -755
rect -539 -765 -535 -755
rect -519 -765 -515 -755
rect -507 -765 -503 -755
rect -499 -765 -495 -755
rect -385 -792 -381 -772
rect -365 -792 -361 -772
rect -348 -776 -344 -766
rect -340 -776 -336 -766
rect -385 -801 -381 -797
rect -375 -801 -371 -797
rect -365 -801 -361 -797
rect -343 -801 -339 -797
rect -605 -868 -601 -858
rect -597 -868 -593 -858
rect -570 -868 -566 -858
rect -550 -868 -546 -858
rect -537 -868 -533 -858
rect -517 -868 -513 -858
rect -505 -868 -501 -858
rect -497 -868 -493 -858
rect -308 -908 -304 -888
rect -288 -908 -280 -888
rect -264 -908 -260 -888
rect -441 -920 -437 -910
rect -433 -920 -429 -910
rect -439 -1062 -435 -1052
rect -431 -1062 -427 -1052
rect -605 -1115 -601 -1105
rect -597 -1115 -593 -1105
rect -570 -1115 -566 -1105
rect -550 -1115 -546 -1105
rect -537 -1115 -533 -1105
rect -517 -1115 -513 -1105
rect -505 -1115 -501 -1105
rect -497 -1115 -493 -1105
rect -384 -1146 -380 -1126
rect -364 -1146 -360 -1126
rect -347 -1130 -343 -1120
rect -339 -1130 -335 -1120
rect -384 -1155 -380 -1151
rect -374 -1155 -370 -1151
rect -364 -1155 -360 -1151
rect -342 -1155 -338 -1151
rect -604 -1225 -600 -1215
rect -596 -1225 -592 -1215
rect -569 -1225 -565 -1215
rect -549 -1225 -545 -1215
rect -536 -1225 -532 -1215
rect -516 -1225 -512 -1215
rect -504 -1225 -500 -1215
rect -496 -1225 -492 -1215
rect -307 -1262 -303 -1242
rect -287 -1262 -279 -1242
rect -263 -1262 -259 -1242
rect -440 -1274 -436 -1264
rect -432 -1274 -428 -1264
rect -81 -1273 -77 -1263
rect -73 -1273 -65 -1263
rect -61 -1273 -57 -1263
rect -44 -1267 -40 -1257
rect -36 -1267 -32 -1257
<< pdcontact >>
rect -441 730 -437 750
rect -433 730 -429 750
rect -603 674 -599 694
rect -583 674 -579 694
rect -568 674 -564 694
rect -560 674 -556 694
rect -535 674 -531 694
rect -527 674 -523 694
rect -503 674 -499 694
rect -495 674 -491 694
rect -384 688 -380 692
rect -376 688 -372 692
rect -368 688 -364 692
rect -349 688 -345 692
rect -386 661 -382 681
rect -378 661 -370 681
rect -366 661 -362 681
rect -349 662 -345 682
rect -341 662 -337 682
rect -605 572 -601 592
rect -585 572 -581 592
rect -570 572 -566 592
rect -562 572 -558 592
rect -537 572 -533 592
rect -529 572 -525 592
rect -505 572 -501 592
rect -497 572 -493 592
rect -309 565 -305 605
rect -289 565 -281 605
rect -265 565 -261 605
rect -442 518 -438 538
rect -434 518 -430 538
rect -441 230 -437 250
rect -433 230 -429 250
rect -603 174 -599 194
rect -583 174 -579 194
rect -568 174 -564 194
rect -560 174 -556 194
rect -535 174 -531 194
rect -527 174 -523 194
rect -503 174 -499 194
rect -495 174 -491 194
rect -384 188 -380 192
rect -376 188 -372 192
rect -368 188 -364 192
rect -349 188 -345 192
rect -386 161 -382 181
rect -378 161 -370 181
rect -366 161 -362 181
rect -349 162 -345 182
rect -341 162 -337 182
rect -605 72 -601 92
rect -585 72 -581 92
rect -570 72 -566 92
rect -562 72 -558 92
rect -537 72 -533 92
rect -529 72 -525 92
rect -505 72 -501 92
rect -497 72 -493 92
rect -309 65 -305 105
rect -289 65 -281 105
rect -265 65 -261 105
rect -442 18 -438 38
rect -434 18 -430 38
rect -442 -217 -438 -197
rect -434 -217 -430 -197
rect -605 -273 -601 -253
rect -585 -273 -581 -253
rect -570 -273 -566 -253
rect -562 -273 -558 -253
rect -537 -273 -533 -253
rect -529 -273 -525 -253
rect -505 -273 -501 -253
rect -497 -273 -493 -253
rect -385 -259 -381 -255
rect -377 -259 -373 -255
rect -369 -259 -365 -255
rect -350 -259 -346 -255
rect -387 -286 -383 -266
rect -379 -286 -371 -266
rect -367 -286 -363 -266
rect -350 -285 -346 -265
rect -342 -285 -338 -265
rect -606 -375 -602 -355
rect -586 -375 -582 -355
rect -571 -375 -567 -355
rect -563 -375 -559 -355
rect -538 -375 -534 -355
rect -530 -375 -526 -355
rect -506 -375 -502 -355
rect -498 -375 -494 -355
rect -310 -382 -306 -342
rect -290 -382 -282 -342
rect -266 -382 -262 -342
rect -443 -429 -439 -409
rect -435 -429 -431 -409
rect -440 -678 -436 -658
rect -432 -678 -428 -658
rect -607 -734 -603 -714
rect -587 -734 -583 -714
rect -572 -734 -568 -714
rect -564 -734 -560 -714
rect -539 -734 -535 -714
rect -531 -734 -527 -714
rect -507 -734 -503 -714
rect -499 -734 -495 -714
rect -383 -720 -379 -716
rect -375 -720 -371 -716
rect -367 -720 -363 -716
rect -348 -720 -344 -716
rect -385 -747 -381 -727
rect -377 -747 -369 -727
rect -365 -747 -361 -727
rect -348 -746 -344 -726
rect -340 -746 -336 -726
rect -605 -837 -601 -817
rect -585 -837 -581 -817
rect -570 -837 -566 -817
rect -562 -837 -558 -817
rect -537 -837 -533 -817
rect -529 -837 -525 -817
rect -505 -837 -501 -817
rect -497 -837 -493 -817
rect -308 -843 -304 -803
rect -288 -843 -280 -803
rect -264 -843 -260 -803
rect -441 -890 -437 -870
rect -433 -890 -429 -870
rect -439 -1032 -435 -1012
rect -431 -1032 -427 -1012
rect -605 -1084 -601 -1064
rect -585 -1084 -581 -1064
rect -570 -1084 -566 -1064
rect -562 -1084 -558 -1064
rect -537 -1084 -533 -1064
rect -529 -1084 -525 -1064
rect -505 -1084 -501 -1064
rect -497 -1084 -493 -1064
rect -382 -1074 -378 -1070
rect -374 -1074 -370 -1070
rect -366 -1074 -362 -1070
rect -347 -1074 -343 -1070
rect -384 -1101 -380 -1081
rect -376 -1101 -368 -1081
rect -364 -1101 -360 -1081
rect -347 -1100 -343 -1080
rect -339 -1100 -335 -1080
rect -604 -1194 -600 -1174
rect -584 -1194 -580 -1174
rect -569 -1194 -565 -1174
rect -561 -1194 -557 -1174
rect -536 -1194 -532 -1174
rect -528 -1194 -524 -1174
rect -504 -1194 -500 -1174
rect -496 -1194 -492 -1174
rect -307 -1197 -303 -1157
rect -287 -1197 -279 -1157
rect -263 -1197 -259 -1157
rect -440 -1244 -436 -1224
rect -432 -1244 -428 -1224
rect -81 -1239 -77 -1199
rect -61 -1239 -57 -1199
rect -44 -1237 -40 -1217
rect -36 -1237 -32 -1217
<< psubstratepcontact >>
rect -603 635 -599 639
rect -568 635 -564 639
rect -559 635 -555 639
rect -548 635 -544 639
rect -535 635 -531 639
rect -525 635 -521 639
rect -515 635 -511 639
rect -503 635 -499 639
rect -605 533 -601 537
rect -570 533 -566 537
rect -561 533 -557 537
rect -550 533 -546 537
rect -537 533 -533 537
rect -527 533 -523 537
rect -517 533 -513 537
rect -505 533 -501 537
rect -309 491 -305 495
rect -299 491 -295 495
rect -287 491 -283 495
rect -275 491 -271 495
rect -265 491 -261 495
rect -603 135 -599 139
rect -568 135 -564 139
rect -559 135 -555 139
rect -548 135 -544 139
rect -535 135 -531 139
rect -525 135 -521 139
rect -515 135 -511 139
rect -503 135 -499 139
rect -605 33 -601 37
rect -570 33 -566 37
rect -561 33 -557 37
rect -550 33 -546 37
rect -537 33 -533 37
rect -527 33 -523 37
rect -517 33 -513 37
rect -505 33 -501 37
rect -309 -9 -305 -5
rect -299 -9 -295 -5
rect -287 -9 -283 -5
rect -275 -9 -271 -5
rect -265 -9 -261 -5
rect -605 -312 -601 -308
rect -570 -312 -566 -308
rect -561 -312 -557 -308
rect -550 -312 -546 -308
rect -537 -312 -533 -308
rect -527 -312 -523 -308
rect -517 -312 -513 -308
rect -505 -312 -501 -308
rect -606 -414 -602 -410
rect -571 -414 -567 -410
rect -562 -414 -558 -410
rect -551 -414 -547 -410
rect -538 -414 -534 -410
rect -528 -414 -524 -410
rect -518 -414 -514 -410
rect -506 -414 -502 -410
rect -310 -456 -306 -452
rect -300 -456 -296 -452
rect -288 -456 -284 -452
rect -276 -456 -272 -452
rect -266 -456 -262 -452
rect -607 -773 -603 -769
rect -572 -773 -568 -769
rect -563 -773 -559 -769
rect -552 -773 -548 -769
rect -539 -773 -535 -769
rect -529 -773 -525 -769
rect -519 -773 -515 -769
rect -507 -773 -503 -769
rect -605 -876 -601 -872
rect -570 -876 -566 -872
rect -561 -876 -557 -872
rect -550 -876 -546 -872
rect -537 -876 -533 -872
rect -527 -876 -523 -872
rect -517 -876 -513 -872
rect -505 -876 -501 -872
rect -308 -917 -304 -913
rect -298 -917 -294 -913
rect -286 -917 -282 -913
rect -274 -917 -270 -913
rect -264 -917 -260 -913
rect -605 -1123 -601 -1119
rect -570 -1123 -566 -1119
rect -561 -1123 -557 -1119
rect -550 -1123 -546 -1119
rect -537 -1123 -533 -1119
rect -527 -1123 -523 -1119
rect -517 -1123 -513 -1119
rect -505 -1123 -501 -1119
rect -604 -1233 -600 -1229
rect -569 -1233 -565 -1229
rect -560 -1233 -556 -1229
rect -549 -1233 -545 -1229
rect -536 -1233 -532 -1229
rect -526 -1233 -522 -1229
rect -516 -1233 -512 -1229
rect -504 -1233 -500 -1229
rect -307 -1271 -303 -1267
rect -297 -1271 -293 -1267
rect -285 -1271 -281 -1267
rect -273 -1271 -269 -1267
rect -263 -1271 -259 -1267
rect -39 -1277 -35 -1273
rect -81 -1283 -77 -1279
rect -71 -1283 -67 -1279
rect -61 -1283 -57 -1279
<< nsubstratencontact >>
rect -603 698 -599 702
rect -593 698 -589 702
rect -583 698 -579 702
rect -563 698 -559 702
rect -535 698 -531 702
rect -503 698 -499 702
rect -309 610 -305 614
rect -299 610 -295 614
rect -287 610 -283 614
rect -276 610 -272 614
rect -265 610 -261 614
rect -605 596 -601 600
rect -595 596 -591 600
rect -585 596 -581 600
rect -565 596 -561 600
rect -537 596 -533 600
rect -505 596 -501 600
rect -603 198 -599 202
rect -593 198 -589 202
rect -583 198 -579 202
rect -563 198 -559 202
rect -535 198 -531 202
rect -503 198 -499 202
rect -309 110 -305 114
rect -299 110 -295 114
rect -287 110 -283 114
rect -276 110 -272 114
rect -265 110 -261 114
rect -605 96 -601 100
rect -595 96 -591 100
rect -585 96 -581 100
rect -565 96 -561 100
rect -537 96 -533 100
rect -505 96 -501 100
rect -605 -249 -601 -245
rect -595 -249 -591 -245
rect -585 -249 -581 -245
rect -565 -249 -561 -245
rect -537 -249 -533 -245
rect -505 -249 -501 -245
rect -310 -337 -306 -333
rect -300 -337 -296 -333
rect -288 -337 -284 -333
rect -277 -337 -273 -333
rect -266 -337 -262 -333
rect -606 -351 -602 -347
rect -596 -351 -592 -347
rect -586 -351 -582 -347
rect -566 -351 -562 -347
rect -538 -351 -534 -347
rect -506 -351 -502 -347
rect -607 -710 -603 -706
rect -597 -710 -593 -706
rect -587 -710 -583 -706
rect -567 -710 -563 -706
rect -539 -710 -535 -706
rect -507 -710 -503 -706
rect -308 -798 -304 -794
rect -298 -798 -294 -794
rect -286 -798 -282 -794
rect -275 -798 -271 -794
rect -264 -798 -260 -794
rect -605 -813 -601 -809
rect -595 -813 -591 -809
rect -585 -813 -581 -809
rect -565 -813 -561 -809
rect -537 -813 -533 -809
rect -505 -813 -501 -809
rect -605 -1060 -601 -1056
rect -595 -1060 -591 -1056
rect -585 -1060 -581 -1056
rect -565 -1060 -561 -1056
rect -537 -1060 -533 -1056
rect -505 -1060 -501 -1056
rect -307 -1152 -303 -1148
rect -297 -1152 -293 -1148
rect -285 -1152 -281 -1148
rect -274 -1152 -270 -1148
rect -263 -1152 -259 -1148
rect -604 -1170 -600 -1166
rect -594 -1170 -590 -1166
rect -584 -1170 -580 -1166
rect -564 -1170 -560 -1166
rect -536 -1170 -532 -1166
rect -504 -1170 -500 -1166
rect -81 -1195 -77 -1191
rect -71 -1195 -67 -1191
rect -61 -1195 -57 -1191
rect -44 -1210 -40 -1206
<< polysilicon >>
rect -436 750 -434 753
rect -436 710 -434 730
rect -598 694 -596 697
rect -586 694 -584 697
rect -563 694 -561 697
rect -530 694 -528 697
rect -498 694 -496 697
rect -436 695 -434 700
rect -381 681 -379 685
rect -369 681 -367 685
rect -344 682 -342 685
rect -598 653 -596 674
rect -598 640 -596 643
rect -586 630 -584 674
rect -563 653 -561 674
rect -551 653 -549 667
rect -530 653 -528 674
rect -518 653 -516 656
rect -498 653 -496 674
rect -563 630 -561 643
rect -551 640 -549 643
rect -530 640 -528 643
rect -518 630 -516 643
rect -498 640 -496 643
rect -381 636 -379 661
rect -369 636 -367 661
rect -344 642 -342 662
rect -586 628 -516 630
rect -344 627 -342 632
rect -381 612 -379 616
rect -369 612 -367 616
rect -304 605 -302 608
rect -292 605 -290 608
rect -280 605 -278 608
rect -268 605 -266 608
rect -600 592 -598 595
rect -588 592 -586 595
rect -565 592 -563 595
rect -532 592 -530 595
rect -500 592 -498 595
rect -600 551 -598 572
rect -600 538 -598 541
rect -588 528 -586 572
rect -565 551 -563 572
rect -553 551 -551 565
rect -532 551 -530 572
rect -520 551 -518 554
rect -500 551 -498 572
rect -304 553 -302 565
rect -292 546 -290 565
rect -280 553 -278 565
rect -268 546 -266 565
rect -565 528 -563 541
rect -553 538 -551 541
rect -532 538 -530 541
rect -520 528 -518 541
rect -500 538 -498 541
rect -437 538 -435 541
rect -588 526 -518 528
rect -304 520 -302 528
rect -292 520 -290 535
rect -280 520 -278 527
rect -268 520 -266 536
rect -437 498 -435 518
rect -304 497 -302 500
rect -292 497 -290 500
rect -280 497 -278 500
rect -268 497 -266 500
rect -437 483 -435 488
rect -436 250 -434 253
rect -436 210 -434 230
rect -598 194 -596 197
rect -586 194 -584 197
rect -563 194 -561 197
rect -530 194 -528 197
rect -498 194 -496 197
rect -436 195 -434 200
rect -381 181 -379 185
rect -369 181 -367 185
rect -344 182 -342 185
rect -598 153 -596 174
rect -598 140 -596 143
rect -586 130 -584 174
rect -563 153 -561 174
rect -551 153 -549 167
rect -530 153 -528 174
rect -518 153 -516 156
rect -498 153 -496 174
rect -563 130 -561 143
rect -551 140 -549 143
rect -530 140 -528 143
rect -518 130 -516 143
rect -498 140 -496 143
rect -381 136 -379 161
rect -369 136 -367 161
rect -344 142 -342 162
rect -586 128 -516 130
rect -344 127 -342 132
rect -381 112 -379 116
rect -369 112 -367 116
rect -304 105 -302 108
rect -292 105 -290 108
rect -280 105 -278 108
rect -268 105 -266 108
rect -600 92 -598 95
rect -588 92 -586 95
rect -565 92 -563 95
rect -532 92 -530 95
rect -500 92 -498 95
rect -600 51 -598 72
rect -600 38 -598 41
rect -588 28 -586 72
rect -565 51 -563 72
rect -553 51 -551 65
rect -532 51 -530 72
rect -520 51 -518 54
rect -500 51 -498 72
rect -304 53 -302 65
rect -292 46 -290 65
rect -280 53 -278 65
rect -268 46 -266 65
rect -565 28 -563 41
rect -553 38 -551 41
rect -532 38 -530 41
rect -520 28 -518 41
rect -500 38 -498 41
rect -437 38 -435 41
rect -588 26 -518 28
rect -304 20 -302 28
rect -292 20 -290 35
rect -280 20 -278 27
rect -268 20 -266 36
rect -437 -2 -435 18
rect -304 -3 -302 0
rect -292 -3 -290 0
rect -280 -3 -278 0
rect -268 -3 -266 0
rect -437 -17 -435 -12
rect -437 -197 -435 -194
rect -437 -237 -435 -217
rect -600 -253 -598 -250
rect -588 -253 -586 -250
rect -565 -253 -563 -250
rect -532 -253 -530 -250
rect -500 -253 -498 -250
rect -437 -252 -435 -247
rect -382 -266 -380 -262
rect -370 -266 -368 -262
rect -345 -265 -343 -262
rect -600 -294 -598 -273
rect -600 -307 -598 -304
rect -588 -317 -586 -273
rect -565 -294 -563 -273
rect -553 -294 -551 -280
rect -532 -294 -530 -273
rect -520 -294 -518 -291
rect -500 -294 -498 -273
rect -565 -317 -563 -304
rect -553 -307 -551 -304
rect -532 -307 -530 -304
rect -520 -317 -518 -304
rect -500 -307 -498 -304
rect -382 -311 -380 -286
rect -370 -311 -368 -286
rect -345 -305 -343 -285
rect -588 -319 -518 -317
rect -345 -320 -343 -315
rect -382 -335 -380 -331
rect -370 -335 -368 -331
rect -305 -342 -303 -339
rect -293 -342 -291 -339
rect -281 -342 -279 -339
rect -269 -342 -267 -339
rect -601 -355 -599 -352
rect -589 -355 -587 -352
rect -566 -355 -564 -352
rect -533 -355 -531 -352
rect -501 -355 -499 -352
rect -601 -396 -599 -375
rect -601 -409 -599 -406
rect -589 -419 -587 -375
rect -566 -396 -564 -375
rect -554 -396 -552 -382
rect -533 -396 -531 -375
rect -521 -396 -519 -393
rect -501 -396 -499 -375
rect -305 -394 -303 -382
rect -293 -401 -291 -382
rect -281 -394 -279 -382
rect -269 -401 -267 -382
rect -566 -419 -564 -406
rect -554 -409 -552 -406
rect -533 -409 -531 -406
rect -521 -419 -519 -406
rect -501 -409 -499 -406
rect -438 -409 -436 -406
rect -589 -421 -519 -419
rect -305 -427 -303 -419
rect -293 -427 -291 -412
rect -281 -427 -279 -420
rect -269 -427 -267 -411
rect -438 -449 -436 -429
rect -305 -450 -303 -447
rect -293 -450 -291 -447
rect -281 -450 -279 -447
rect -269 -450 -267 -447
rect -438 -464 -436 -459
rect -435 -658 -433 -655
rect -435 -698 -433 -678
rect -602 -714 -600 -711
rect -590 -714 -588 -711
rect -567 -714 -565 -711
rect -534 -714 -532 -711
rect -502 -714 -500 -711
rect -435 -713 -433 -708
rect -380 -727 -378 -723
rect -368 -727 -366 -723
rect -343 -726 -341 -723
rect -602 -755 -600 -734
rect -602 -768 -600 -765
rect -590 -778 -588 -734
rect -567 -755 -565 -734
rect -555 -755 -553 -741
rect -534 -755 -532 -734
rect -522 -755 -520 -752
rect -502 -755 -500 -734
rect -567 -778 -565 -765
rect -555 -768 -553 -765
rect -534 -768 -532 -765
rect -522 -778 -520 -765
rect -502 -768 -500 -765
rect -380 -772 -378 -747
rect -368 -772 -366 -747
rect -343 -766 -341 -746
rect -590 -780 -520 -778
rect -343 -781 -341 -776
rect -380 -796 -378 -792
rect -368 -796 -366 -792
rect -303 -803 -301 -800
rect -291 -803 -289 -800
rect -279 -803 -277 -800
rect -267 -803 -265 -800
rect -600 -817 -598 -814
rect -588 -817 -586 -814
rect -565 -817 -563 -814
rect -532 -817 -530 -814
rect -500 -817 -498 -814
rect -600 -858 -598 -837
rect -600 -871 -598 -868
rect -588 -881 -586 -837
rect -565 -858 -563 -837
rect -553 -858 -551 -844
rect -532 -858 -530 -837
rect -520 -858 -518 -855
rect -500 -858 -498 -837
rect -303 -855 -301 -843
rect -291 -862 -289 -843
rect -279 -855 -277 -843
rect -267 -862 -265 -843
rect -565 -881 -563 -868
rect -553 -871 -551 -868
rect -532 -871 -530 -868
rect -520 -881 -518 -868
rect -500 -871 -498 -868
rect -436 -870 -434 -867
rect -588 -883 -518 -881
rect -303 -888 -301 -880
rect -291 -888 -289 -873
rect -279 -888 -277 -881
rect -267 -888 -265 -872
rect -436 -910 -434 -890
rect -303 -911 -301 -908
rect -291 -911 -289 -908
rect -279 -911 -277 -908
rect -267 -911 -265 -908
rect -436 -925 -434 -920
rect -434 -1012 -432 -1009
rect -434 -1052 -432 -1032
rect -600 -1064 -598 -1061
rect -588 -1064 -586 -1061
rect -565 -1064 -563 -1061
rect -532 -1064 -530 -1061
rect -500 -1064 -498 -1061
rect -434 -1067 -432 -1062
rect -379 -1081 -377 -1077
rect -367 -1081 -365 -1077
rect -342 -1080 -340 -1077
rect -600 -1105 -598 -1084
rect -600 -1118 -598 -1115
rect -588 -1128 -586 -1084
rect -565 -1105 -563 -1084
rect -553 -1105 -551 -1091
rect -532 -1105 -530 -1084
rect -520 -1105 -518 -1102
rect -500 -1105 -498 -1084
rect -565 -1128 -563 -1115
rect -553 -1118 -551 -1115
rect -532 -1118 -530 -1115
rect -520 -1128 -518 -1115
rect -500 -1118 -498 -1115
rect -379 -1126 -377 -1101
rect -367 -1126 -365 -1101
rect -342 -1120 -340 -1100
rect -588 -1130 -518 -1128
rect -342 -1135 -340 -1130
rect -379 -1150 -377 -1146
rect -367 -1150 -365 -1146
rect -302 -1157 -300 -1154
rect -290 -1157 -288 -1154
rect -278 -1157 -276 -1154
rect -266 -1157 -264 -1154
rect -599 -1174 -597 -1171
rect -587 -1174 -585 -1171
rect -564 -1174 -562 -1171
rect -531 -1174 -529 -1171
rect -499 -1174 -497 -1171
rect -599 -1215 -597 -1194
rect -599 -1228 -597 -1225
rect -587 -1238 -585 -1194
rect -564 -1215 -562 -1194
rect -552 -1215 -550 -1201
rect -531 -1215 -529 -1194
rect -519 -1215 -517 -1212
rect -499 -1215 -497 -1194
rect -302 -1209 -300 -1197
rect -290 -1216 -288 -1197
rect -278 -1209 -276 -1197
rect -266 -1216 -264 -1197
rect -76 -1199 -74 -1196
rect -64 -1199 -62 -1196
rect -435 -1224 -433 -1221
rect -564 -1238 -562 -1225
rect -552 -1228 -550 -1225
rect -531 -1228 -529 -1225
rect -519 -1238 -517 -1225
rect -499 -1228 -497 -1225
rect -587 -1240 -517 -1238
rect -302 -1242 -300 -1234
rect -290 -1242 -288 -1227
rect -278 -1242 -276 -1235
rect -266 -1242 -264 -1226
rect -39 -1217 -37 -1214
rect -435 -1264 -433 -1244
rect -302 -1265 -300 -1262
rect -290 -1265 -288 -1262
rect -278 -1265 -276 -1262
rect -266 -1265 -264 -1262
rect -76 -1263 -74 -1239
rect -64 -1263 -62 -1239
rect -39 -1257 -37 -1237
rect -39 -1272 -37 -1267
rect -435 -1279 -433 -1274
rect -76 -1276 -74 -1273
rect -64 -1276 -62 -1273
<< polycontact >>
rect -440 715 -436 719
rect -602 656 -598 660
rect -590 663 -586 667
rect -555 662 -551 666
rect -534 662 -530 666
rect -502 662 -498 666
rect -386 649 -381 653
rect -375 640 -369 644
rect -348 647 -344 651
rect -604 554 -600 558
rect -592 561 -588 565
rect -557 560 -553 564
rect -536 560 -532 564
rect -504 560 -500 564
rect -308 554 -304 558
rect -296 547 -292 551
rect -278 554 -274 558
rect -266 547 -262 551
rect -296 530 -292 534
rect -308 523 -304 527
rect -278 523 -274 527
rect -266 530 -262 534
rect -441 503 -437 507
rect -440 215 -436 219
rect -602 156 -598 160
rect -590 163 -586 167
rect -555 162 -551 166
rect -534 162 -530 166
rect -502 162 -498 166
rect -386 149 -381 153
rect -375 140 -369 144
rect -348 147 -344 151
rect -604 54 -600 58
rect -592 61 -588 65
rect -557 60 -553 64
rect -536 60 -532 64
rect -504 60 -500 64
rect -308 54 -304 58
rect -296 47 -292 51
rect -278 54 -274 58
rect -266 47 -262 51
rect -296 30 -292 34
rect -308 23 -304 27
rect -278 23 -274 27
rect -266 30 -262 34
rect -441 3 -437 7
rect -441 -232 -437 -228
rect -604 -291 -600 -287
rect -592 -284 -588 -280
rect -557 -285 -553 -281
rect -536 -285 -532 -281
rect -504 -285 -500 -281
rect -387 -298 -382 -294
rect -376 -307 -370 -303
rect -349 -300 -345 -296
rect -605 -393 -601 -389
rect -593 -386 -589 -382
rect -558 -387 -554 -383
rect -537 -387 -533 -383
rect -505 -387 -501 -383
rect -309 -393 -305 -389
rect -297 -400 -293 -396
rect -279 -393 -275 -389
rect -267 -400 -263 -396
rect -297 -417 -293 -413
rect -309 -424 -305 -420
rect -279 -424 -275 -420
rect -267 -417 -263 -413
rect -442 -444 -438 -440
rect -439 -693 -435 -689
rect -606 -752 -602 -748
rect -594 -745 -590 -741
rect -559 -746 -555 -742
rect -538 -746 -534 -742
rect -506 -746 -502 -742
rect -385 -759 -380 -755
rect -374 -768 -368 -764
rect -347 -761 -343 -757
rect -604 -855 -600 -851
rect -592 -848 -588 -844
rect -557 -849 -553 -845
rect -536 -849 -532 -845
rect -504 -849 -500 -845
rect -307 -854 -303 -850
rect -295 -861 -291 -857
rect -277 -854 -273 -850
rect -265 -861 -261 -857
rect -295 -878 -291 -874
rect -307 -885 -303 -881
rect -277 -885 -273 -881
rect -265 -878 -261 -874
rect -440 -905 -436 -901
rect -438 -1047 -434 -1043
rect -604 -1102 -600 -1098
rect -592 -1095 -588 -1091
rect -557 -1096 -553 -1092
rect -536 -1096 -532 -1092
rect -504 -1096 -500 -1092
rect -384 -1113 -379 -1109
rect -373 -1122 -367 -1118
rect -346 -1115 -342 -1111
rect -603 -1212 -599 -1208
rect -591 -1205 -587 -1201
rect -556 -1206 -552 -1202
rect -535 -1206 -531 -1202
rect -503 -1206 -499 -1202
rect -306 -1208 -302 -1204
rect -294 -1215 -290 -1211
rect -276 -1208 -272 -1204
rect -264 -1215 -260 -1211
rect -294 -1232 -290 -1228
rect -306 -1239 -302 -1235
rect -276 -1239 -272 -1235
rect -264 -1232 -260 -1228
rect -439 -1259 -435 -1255
rect -81 -1260 -76 -1256
rect -69 -1253 -64 -1249
rect -43 -1252 -39 -1248
<< metal1 >>
rect -638 667 -634 785
rect -448 756 -422 761
rect -441 750 -437 756
rect -433 719 -429 730
rect -475 715 -440 719
rect -433 715 -232 719
rect -599 698 -593 702
rect -589 698 -583 702
rect -579 698 -563 702
rect -559 698 -535 702
rect -531 698 -503 702
rect -499 698 -485 702
rect -603 694 -599 698
rect -568 694 -564 698
rect -535 694 -531 698
rect -503 694 -499 698
rect -556 674 -544 694
rect -523 674 -511 694
rect -638 663 -590 667
rect -583 666 -579 674
rect -548 666 -544 674
rect -515 666 -511 674
rect -495 666 -491 674
rect -475 666 -470 715
rect -433 710 -429 715
rect -441 694 -437 700
rect -441 690 -429 694
rect -386 692 -330 694
rect -638 565 -634 663
rect -583 662 -555 666
rect -548 662 -534 666
rect -515 662 -502 666
rect -495 662 -470 666
rect -609 656 -602 660
rect -583 653 -579 662
rect -548 653 -544 662
rect -515 653 -511 662
rect -495 653 -491 662
rect -591 643 -579 653
rect -475 656 -470 662
rect -386 688 -384 692
rect -380 688 -376 692
rect -372 688 -368 692
rect -364 688 -349 692
rect -345 688 -330 692
rect -386 686 -362 688
rect -386 681 -382 686
rect -366 681 -362 686
rect -349 682 -345 688
rect -475 649 -439 656
rect -432 653 -427 656
rect -378 654 -370 661
rect -432 649 -386 653
rect -378 651 -362 654
rect -341 651 -337 662
rect -378 650 -348 651
rect -366 647 -348 650
rect -341 647 -326 651
rect -603 639 -599 643
rect -568 639 -564 643
rect -535 639 -531 643
rect -503 639 -499 643
rect -474 640 -375 644
rect -599 635 -568 639
rect -564 635 -559 639
rect -555 635 -548 639
rect -544 635 -535 639
rect -531 635 -525 639
rect -521 635 -515 639
rect -511 635 -503 639
rect -499 635 -491 639
rect -601 596 -595 600
rect -591 596 -585 600
rect -581 596 -565 600
rect -561 596 -537 600
rect -533 596 -505 600
rect -501 596 -487 600
rect -605 592 -601 596
rect -570 592 -566 596
rect -537 592 -533 596
rect -505 592 -501 596
rect -558 572 -546 592
rect -525 572 -513 592
rect -638 561 -592 565
rect -585 564 -581 572
rect -550 564 -546 572
rect -517 564 -513 572
rect -497 564 -493 572
rect -474 588 -470 640
rect -366 636 -362 647
rect -341 642 -337 647
rect -349 626 -345 632
rect -386 611 -382 616
rect -349 611 -336 626
rect -392 607 -386 611
rect -382 607 -376 611
rect -372 607 -366 611
rect -362 607 -344 611
rect -340 607 -336 611
rect -326 621 -248 626
rect -326 588 -322 621
rect -474 584 -322 588
rect -305 610 -299 614
rect -295 610 -287 614
rect -283 610 -276 614
rect -272 610 -265 614
rect -309 609 -261 610
rect -309 605 -305 609
rect -265 605 -261 609
rect -474 564 -470 584
rect -638 167 -634 561
rect -585 560 -557 564
rect -550 560 -536 564
rect -517 560 -504 564
rect -497 560 -470 564
rect -611 554 -604 558
rect -585 551 -581 560
rect -550 551 -546 560
rect -517 551 -513 560
rect -497 551 -493 560
rect -593 541 -581 551
rect -605 537 -601 541
rect -570 537 -566 541
rect -537 537 -533 541
rect -505 537 -501 541
rect -601 533 -570 537
rect -566 533 -561 537
rect -557 533 -550 537
rect -546 533 -537 537
rect -533 533 -527 537
rect -523 533 -517 537
rect -513 533 -505 537
rect -501 533 -493 537
rect -475 507 -470 560
rect -432 555 -308 558
rect -449 544 -423 549
rect -442 538 -438 544
rect -340 534 -336 555
rect -320 554 -308 555
rect -308 547 -296 551
rect -289 543 -281 565
rect -252 558 -248 621
rect -274 554 -248 558
rect -236 554 -232 715
rect -262 547 -242 551
rect -234 547 -232 554
rect -210 666 -175 670
rect -210 589 -206 666
rect -179 655 -175 661
rect -210 585 -175 589
rect -210 543 -206 585
rect -289 539 -205 543
rect -289 538 -213 539
rect -340 530 -296 534
rect -434 507 -430 518
rect -328 523 -308 527
rect -475 503 -441 507
rect -434 503 -363 507
rect -475 468 -470 503
rect -434 498 -430 503
rect -442 482 -438 488
rect -442 478 -430 482
rect -328 468 -323 523
rect -289 520 -281 538
rect -262 530 -242 534
rect -274 523 -252 527
rect -309 496 -305 500
rect -265 496 -261 500
rect -309 495 -261 496
rect -305 491 -299 495
rect -295 491 -287 495
rect -283 491 -275 495
rect -271 491 -265 495
rect -475 464 -323 468
rect -255 457 -252 523
rect -352 448 -239 457
rect -448 256 -422 261
rect -441 250 -437 256
rect -433 219 -429 230
rect -475 215 -440 219
rect -433 215 -232 219
rect -599 198 -593 202
rect -589 198 -583 202
rect -579 198 -563 202
rect -559 198 -535 202
rect -531 198 -503 202
rect -499 198 -485 202
rect -603 194 -599 198
rect -568 194 -564 198
rect -535 194 -531 198
rect -503 194 -499 198
rect -556 174 -544 194
rect -523 174 -511 194
rect -638 163 -590 167
rect -583 166 -579 174
rect -548 166 -544 174
rect -515 166 -511 174
rect -495 166 -491 174
rect -475 166 -470 215
rect -433 210 -429 215
rect -441 194 -437 200
rect -441 190 -429 194
rect -386 192 -330 194
rect -638 65 -634 163
rect -583 162 -555 166
rect -548 162 -534 166
rect -515 162 -502 166
rect -495 162 -470 166
rect -609 156 -602 160
rect -583 153 -579 162
rect -548 153 -544 162
rect -515 153 -511 162
rect -495 153 -491 162
rect -591 143 -579 153
rect -475 156 -470 162
rect -386 188 -384 192
rect -380 188 -376 192
rect -372 188 -368 192
rect -364 188 -349 192
rect -345 188 -330 192
rect -386 186 -362 188
rect -386 181 -382 186
rect -366 181 -362 186
rect -349 182 -345 188
rect -475 149 -439 156
rect -432 153 -427 156
rect -378 154 -370 161
rect -432 149 -386 153
rect -378 151 -362 154
rect -341 151 -337 162
rect -378 150 -348 151
rect -366 147 -348 150
rect -341 147 -326 151
rect -603 139 -599 143
rect -568 139 -564 143
rect -535 139 -531 143
rect -503 139 -499 143
rect -474 140 -375 144
rect -599 135 -568 139
rect -564 135 -559 139
rect -555 135 -548 139
rect -544 135 -535 139
rect -531 135 -525 139
rect -521 135 -515 139
rect -511 135 -503 139
rect -499 135 -491 139
rect -601 96 -595 100
rect -591 96 -585 100
rect -581 96 -565 100
rect -561 96 -537 100
rect -533 96 -505 100
rect -501 96 -487 100
rect -605 92 -601 96
rect -570 92 -566 96
rect -537 92 -533 96
rect -505 92 -501 96
rect -558 72 -546 92
rect -525 72 -513 92
rect -638 61 -592 65
rect -585 64 -581 72
rect -550 64 -546 72
rect -517 64 -513 72
rect -497 64 -493 72
rect -474 88 -470 140
rect -366 136 -362 147
rect -341 142 -337 147
rect -349 126 -345 132
rect -386 111 -382 116
rect -349 111 -336 126
rect -392 107 -386 111
rect -382 107 -376 111
rect -372 107 -366 111
rect -362 107 -344 111
rect -340 107 -336 111
rect -326 121 -248 126
rect -326 88 -322 121
rect -474 84 -322 88
rect -305 110 -299 114
rect -295 110 -287 114
rect -283 110 -276 114
rect -272 110 -265 114
rect -309 109 -261 110
rect -309 105 -305 109
rect -265 105 -261 109
rect -474 64 -470 84
rect -638 -280 -634 61
rect -585 60 -557 64
rect -550 60 -536 64
rect -517 60 -504 64
rect -497 60 -470 64
rect -611 54 -604 58
rect -585 51 -581 60
rect -550 51 -546 60
rect -517 51 -513 60
rect -497 51 -493 60
rect -593 41 -581 51
rect -605 37 -601 41
rect -570 37 -566 41
rect -537 37 -533 41
rect -505 37 -501 41
rect -601 33 -570 37
rect -566 33 -561 37
rect -557 33 -550 37
rect -546 33 -537 37
rect -533 33 -527 37
rect -523 33 -517 37
rect -513 33 -505 37
rect -501 33 -493 37
rect -475 7 -470 60
rect -432 55 -308 58
rect -449 44 -423 49
rect -442 38 -438 44
rect -340 34 -336 55
rect -320 54 -308 55
rect -308 47 -296 51
rect -289 43 -281 65
rect -252 58 -248 121
rect -274 54 -248 58
rect -236 54 -232 215
rect -262 47 -242 51
rect -234 47 -232 54
rect -210 166 -175 170
rect -210 89 -206 166
rect -179 155 -175 161
rect -210 85 -175 89
rect -210 43 -206 85
rect -289 39 -205 43
rect -289 38 -213 39
rect -340 30 -296 34
rect -434 7 -430 18
rect -328 23 -308 27
rect -475 3 -441 7
rect -434 3 -363 7
rect -475 -32 -470 3
rect -434 -2 -430 3
rect -442 -18 -438 -12
rect -442 -22 -430 -18
rect -328 -32 -323 23
rect -289 20 -281 38
rect -262 30 -242 34
rect -274 23 -252 27
rect -309 -4 -305 0
rect -265 -4 -261 0
rect -309 -5 -261 -4
rect -305 -9 -299 -5
rect -295 -9 -287 -5
rect -283 -9 -275 -5
rect -271 -9 -265 -5
rect -475 -36 -323 -32
rect -255 -43 -252 23
rect -352 -52 -239 -43
rect -449 -191 -423 -186
rect -442 -197 -438 -191
rect -434 -228 -430 -217
rect -476 -232 -441 -228
rect -434 -232 -233 -228
rect -601 -249 -595 -245
rect -591 -249 -585 -245
rect -581 -249 -565 -245
rect -561 -249 -537 -245
rect -533 -249 -505 -245
rect -501 -249 -487 -245
rect -605 -253 -601 -249
rect -570 -253 -566 -249
rect -537 -253 -533 -249
rect -505 -253 -501 -249
rect -558 -273 -546 -253
rect -525 -273 -513 -253
rect -638 -284 -592 -280
rect -585 -281 -581 -273
rect -550 -281 -546 -273
rect -517 -281 -513 -273
rect -497 -281 -493 -273
rect -476 -281 -471 -232
rect -434 -237 -430 -232
rect -442 -253 -438 -247
rect -442 -257 -430 -253
rect -387 -255 -331 -253
rect -638 -382 -634 -284
rect -585 -285 -557 -281
rect -550 -285 -536 -281
rect -517 -285 -504 -281
rect -497 -285 -471 -281
rect -611 -291 -604 -287
rect -585 -294 -581 -285
rect -550 -294 -546 -285
rect -517 -294 -513 -285
rect -497 -294 -493 -285
rect -593 -304 -581 -294
rect -476 -291 -471 -285
rect -387 -259 -385 -255
rect -381 -259 -377 -255
rect -373 -259 -369 -255
rect -365 -259 -350 -255
rect -346 -259 -331 -255
rect -387 -261 -363 -259
rect -387 -266 -383 -261
rect -367 -266 -363 -261
rect -350 -265 -346 -259
rect -476 -298 -440 -291
rect -433 -294 -428 -291
rect -379 -293 -371 -286
rect -433 -298 -387 -294
rect -379 -296 -363 -293
rect -342 -296 -338 -285
rect -379 -297 -349 -296
rect -367 -300 -349 -297
rect -342 -300 -312 -296
rect -605 -308 -601 -304
rect -570 -308 -566 -304
rect -537 -308 -533 -304
rect -505 -308 -501 -304
rect -475 -307 -376 -303
rect -601 -312 -570 -308
rect -566 -312 -561 -308
rect -557 -312 -550 -308
rect -546 -312 -537 -308
rect -533 -312 -527 -308
rect -523 -312 -517 -308
rect -513 -312 -505 -308
rect -501 -312 -493 -308
rect -602 -351 -596 -347
rect -592 -351 -586 -347
rect -582 -351 -566 -347
rect -562 -351 -538 -347
rect -534 -351 -506 -347
rect -502 -351 -488 -347
rect -606 -355 -602 -351
rect -571 -355 -567 -351
rect -538 -355 -534 -351
rect -506 -355 -502 -351
rect -559 -375 -547 -355
rect -526 -375 -514 -355
rect -638 -386 -593 -382
rect -586 -383 -582 -375
rect -551 -383 -547 -375
rect -518 -383 -514 -375
rect -498 -383 -494 -375
rect -475 -359 -471 -307
rect -367 -311 -363 -300
rect -342 -305 -338 -300
rect -350 -321 -346 -315
rect -387 -336 -383 -331
rect -350 -336 -337 -321
rect -393 -340 -387 -336
rect -383 -340 -377 -336
rect -373 -340 -367 -336
rect -363 -340 -345 -336
rect -341 -340 -337 -336
rect -327 -326 -249 -321
rect -327 -359 -323 -326
rect -475 -363 -323 -359
rect -306 -337 -300 -333
rect -296 -337 -288 -333
rect -284 -337 -277 -333
rect -273 -337 -266 -333
rect -310 -338 -262 -337
rect -310 -342 -306 -338
rect -266 -342 -262 -338
rect -475 -383 -471 -363
rect -638 -741 -634 -386
rect -586 -387 -558 -383
rect -551 -387 -537 -383
rect -518 -387 -505 -383
rect -498 -387 -471 -383
rect -612 -393 -605 -389
rect -586 -396 -582 -387
rect -551 -396 -547 -387
rect -518 -396 -514 -387
rect -498 -396 -494 -387
rect -594 -406 -582 -396
rect -606 -410 -602 -406
rect -571 -410 -567 -406
rect -538 -410 -534 -406
rect -506 -410 -502 -406
rect -602 -414 -571 -410
rect -567 -414 -562 -410
rect -558 -414 -551 -410
rect -547 -414 -538 -410
rect -534 -414 -528 -410
rect -524 -414 -518 -410
rect -514 -414 -506 -410
rect -502 -414 -494 -410
rect -476 -440 -471 -387
rect -433 -392 -309 -389
rect -450 -403 -424 -398
rect -443 -409 -439 -403
rect -341 -413 -337 -392
rect -321 -393 -309 -392
rect -309 -400 -297 -396
rect -290 -404 -282 -382
rect -253 -389 -249 -326
rect -275 -393 -249 -389
rect -237 -393 -233 -232
rect -263 -400 -243 -396
rect -235 -400 -233 -393
rect -187 -279 -175 -275
rect -187 -347 -182 -279
rect -187 -351 -175 -347
rect -187 -404 -182 -351
rect -290 -409 -182 -404
rect -341 -417 -297 -413
rect -435 -440 -431 -429
rect -329 -424 -309 -420
rect -476 -444 -442 -440
rect -435 -444 -364 -440
rect -476 -479 -471 -444
rect -435 -449 -431 -444
rect -443 -465 -439 -459
rect -443 -469 -431 -465
rect -329 -479 -324 -424
rect -290 -427 -282 -409
rect -263 -417 -243 -413
rect -275 -424 -253 -420
rect -310 -451 -306 -447
rect -266 -451 -262 -447
rect -310 -452 -262 -451
rect -306 -456 -300 -452
rect -296 -456 -288 -452
rect -284 -456 -276 -452
rect -272 -456 -266 -452
rect -476 -483 -324 -479
rect -256 -490 -253 -424
rect -353 -499 -240 -490
rect -447 -652 -421 -647
rect -440 -658 -436 -652
rect -432 -689 -428 -678
rect -474 -693 -439 -689
rect -432 -693 -231 -689
rect -603 -710 -597 -706
rect -593 -710 -587 -706
rect -583 -710 -567 -706
rect -563 -710 -539 -706
rect -535 -710 -507 -706
rect -503 -710 -489 -706
rect -607 -714 -603 -710
rect -572 -714 -568 -710
rect -539 -714 -535 -710
rect -507 -714 -503 -710
rect -560 -734 -548 -714
rect -527 -734 -515 -714
rect -638 -745 -594 -741
rect -587 -742 -583 -734
rect -552 -742 -548 -734
rect -519 -742 -515 -734
rect -499 -742 -495 -734
rect -474 -742 -469 -693
rect -432 -698 -428 -693
rect -440 -714 -436 -708
rect -440 -718 -428 -714
rect -385 -716 -329 -714
rect -638 -844 -634 -745
rect -587 -746 -559 -742
rect -552 -746 -538 -742
rect -519 -746 -506 -742
rect -499 -746 -469 -742
rect -613 -752 -606 -748
rect -587 -755 -583 -746
rect -552 -755 -548 -746
rect -519 -755 -515 -746
rect -499 -755 -495 -746
rect -595 -765 -583 -755
rect -474 -752 -469 -746
rect -385 -720 -383 -716
rect -379 -720 -375 -716
rect -371 -720 -367 -716
rect -363 -720 -348 -716
rect -344 -720 -329 -716
rect -385 -722 -361 -720
rect -385 -727 -381 -722
rect -365 -727 -361 -722
rect -348 -726 -344 -720
rect -474 -759 -438 -752
rect -431 -755 -426 -752
rect -377 -754 -369 -747
rect -431 -759 -385 -755
rect -377 -757 -361 -754
rect -340 -757 -336 -746
rect -377 -758 -347 -757
rect -365 -761 -347 -758
rect -340 -761 -317 -757
rect -607 -769 -603 -765
rect -572 -769 -568 -765
rect -539 -769 -535 -765
rect -507 -769 -503 -765
rect -473 -768 -374 -764
rect -603 -773 -572 -769
rect -568 -773 -563 -769
rect -559 -773 -552 -769
rect -548 -773 -539 -769
rect -535 -773 -529 -769
rect -525 -773 -519 -769
rect -515 -773 -507 -769
rect -503 -773 -495 -769
rect -601 -813 -595 -809
rect -591 -813 -585 -809
rect -581 -813 -565 -809
rect -561 -813 -537 -809
rect -533 -813 -505 -809
rect -501 -813 -487 -809
rect -605 -817 -601 -813
rect -570 -817 -566 -813
rect -537 -817 -533 -813
rect -505 -817 -501 -813
rect -558 -837 -546 -817
rect -525 -837 -513 -817
rect -638 -848 -592 -844
rect -585 -845 -581 -837
rect -550 -845 -546 -837
rect -517 -845 -513 -837
rect -497 -845 -493 -837
rect -473 -820 -469 -768
rect -365 -772 -361 -761
rect -340 -766 -336 -761
rect -348 -782 -344 -776
rect -385 -797 -381 -792
rect -348 -797 -335 -782
rect -391 -801 -385 -797
rect -381 -801 -375 -797
rect -371 -801 -365 -797
rect -361 -801 -343 -797
rect -339 -801 -335 -797
rect -325 -787 -247 -782
rect -325 -820 -321 -787
rect -473 -824 -321 -820
rect -304 -798 -298 -794
rect -294 -798 -286 -794
rect -282 -798 -275 -794
rect -271 -798 -264 -794
rect -308 -799 -260 -798
rect -308 -803 -304 -799
rect -264 -803 -260 -799
rect -473 -845 -469 -824
rect -638 -980 -634 -848
rect -585 -849 -557 -845
rect -550 -849 -536 -845
rect -517 -849 -504 -845
rect -497 -849 -469 -845
rect -611 -855 -604 -851
rect -585 -858 -581 -849
rect -550 -858 -546 -849
rect -517 -858 -513 -849
rect -497 -858 -493 -849
rect -593 -868 -581 -858
rect -605 -872 -601 -868
rect -570 -872 -566 -868
rect -537 -872 -533 -868
rect -505 -872 -501 -868
rect -601 -876 -570 -872
rect -566 -876 -561 -872
rect -557 -876 -550 -872
rect -546 -876 -537 -872
rect -533 -876 -527 -872
rect -523 -876 -517 -872
rect -513 -876 -505 -872
rect -501 -876 -493 -872
rect -474 -901 -469 -849
rect -431 -853 -307 -850
rect -448 -864 -422 -859
rect -441 -870 -437 -864
rect -339 -874 -335 -853
rect -319 -854 -307 -853
rect -307 -861 -295 -857
rect -288 -865 -280 -843
rect -251 -850 -247 -787
rect -273 -854 -247 -850
rect -235 -854 -231 -693
rect -261 -861 -241 -857
rect -233 -861 -231 -854
rect -288 -870 -175 -865
rect -339 -878 -295 -874
rect -433 -901 -429 -890
rect -327 -885 -307 -881
rect -474 -905 -440 -901
rect -433 -905 -362 -901
rect -474 -940 -469 -905
rect -433 -910 -429 -905
rect -441 -926 -437 -920
rect -441 -930 -429 -926
rect -327 -940 -322 -885
rect -288 -888 -280 -870
rect -261 -878 -241 -874
rect -273 -885 -251 -881
rect -308 -912 -304 -908
rect -264 -912 -260 -908
rect -308 -913 -260 -912
rect -304 -917 -298 -913
rect -294 -917 -286 -913
rect -282 -917 -274 -913
rect -270 -917 -264 -913
rect -474 -944 -322 -940
rect -254 -951 -251 -885
rect -351 -960 -238 -951
rect -715 -984 -634 -980
rect -715 -1043 -711 -984
rect -446 -1006 -420 -1001
rect -439 -1012 -435 -1006
rect -431 -1043 -427 -1032
rect -715 -1047 -623 -1043
rect -627 -1091 -623 -1047
rect -473 -1047 -438 -1043
rect -431 -1047 -230 -1043
rect -601 -1060 -595 -1056
rect -591 -1060 -585 -1056
rect -581 -1060 -565 -1056
rect -561 -1060 -537 -1056
rect -533 -1060 -505 -1056
rect -501 -1060 -487 -1056
rect -605 -1064 -601 -1060
rect -570 -1064 -566 -1060
rect -537 -1064 -533 -1060
rect -505 -1064 -501 -1060
rect -558 -1084 -546 -1064
rect -525 -1084 -513 -1064
rect -627 -1095 -592 -1091
rect -585 -1092 -581 -1084
rect -550 -1092 -546 -1084
rect -517 -1092 -513 -1084
rect -497 -1092 -493 -1084
rect -473 -1092 -468 -1047
rect -431 -1052 -427 -1047
rect -439 -1068 -435 -1062
rect -439 -1072 -427 -1068
rect -384 -1070 -328 -1068
rect -627 -1201 -623 -1095
rect -585 -1096 -557 -1092
rect -550 -1096 -536 -1092
rect -517 -1096 -504 -1092
rect -497 -1096 -468 -1092
rect -611 -1102 -604 -1098
rect -585 -1105 -581 -1096
rect -550 -1105 -546 -1096
rect -517 -1105 -513 -1096
rect -497 -1105 -493 -1096
rect -593 -1115 -581 -1105
rect -473 -1106 -468 -1096
rect -384 -1074 -382 -1070
rect -378 -1074 -374 -1070
rect -370 -1074 -366 -1070
rect -362 -1074 -347 -1070
rect -343 -1074 -328 -1070
rect -384 -1076 -360 -1074
rect -384 -1081 -380 -1076
rect -364 -1081 -360 -1076
rect -347 -1080 -343 -1074
rect -473 -1113 -437 -1106
rect -430 -1109 -425 -1106
rect -376 -1108 -368 -1101
rect -430 -1113 -384 -1109
rect -376 -1111 -360 -1108
rect -339 -1111 -335 -1100
rect -376 -1112 -346 -1111
rect -364 -1115 -346 -1112
rect -339 -1115 -322 -1111
rect -605 -1119 -601 -1115
rect -570 -1119 -566 -1115
rect -537 -1119 -533 -1115
rect -505 -1119 -501 -1115
rect -601 -1123 -570 -1119
rect -566 -1123 -561 -1119
rect -557 -1123 -550 -1119
rect -546 -1123 -537 -1119
rect -533 -1123 -527 -1119
rect -523 -1123 -517 -1119
rect -513 -1123 -505 -1119
rect -501 -1123 -493 -1119
rect -472 -1122 -373 -1118
rect -600 -1170 -594 -1166
rect -590 -1170 -584 -1166
rect -580 -1170 -564 -1166
rect -560 -1170 -536 -1166
rect -532 -1170 -504 -1166
rect -500 -1170 -486 -1166
rect -604 -1174 -600 -1170
rect -569 -1174 -565 -1170
rect -536 -1174 -532 -1170
rect -504 -1174 -500 -1170
rect -472 -1174 -468 -1122
rect -364 -1126 -360 -1115
rect -339 -1120 -335 -1115
rect -347 -1136 -343 -1130
rect -384 -1151 -380 -1146
rect -347 -1151 -334 -1136
rect -390 -1155 -384 -1151
rect -380 -1155 -374 -1151
rect -370 -1155 -364 -1151
rect -360 -1155 -342 -1151
rect -338 -1155 -334 -1151
rect -324 -1141 -246 -1136
rect -324 -1174 -320 -1141
rect -557 -1194 -545 -1174
rect -524 -1194 -512 -1174
rect -627 -1205 -591 -1201
rect -584 -1202 -580 -1194
rect -549 -1202 -545 -1194
rect -516 -1202 -512 -1194
rect -496 -1202 -492 -1194
rect -472 -1178 -320 -1174
rect -303 -1152 -297 -1148
rect -293 -1152 -285 -1148
rect -281 -1152 -274 -1148
rect -270 -1152 -263 -1148
rect -307 -1153 -259 -1152
rect -307 -1157 -303 -1153
rect -263 -1157 -259 -1153
rect -472 -1202 -468 -1178
rect -584 -1206 -556 -1202
rect -549 -1206 -535 -1202
rect -516 -1206 -503 -1202
rect -496 -1206 -468 -1202
rect -610 -1212 -603 -1208
rect -584 -1215 -580 -1206
rect -549 -1215 -545 -1206
rect -516 -1215 -512 -1206
rect -496 -1215 -492 -1206
rect -592 -1225 -580 -1215
rect -604 -1229 -600 -1225
rect -569 -1229 -565 -1225
rect -536 -1229 -532 -1225
rect -504 -1229 -500 -1225
rect -600 -1233 -569 -1229
rect -565 -1233 -560 -1229
rect -556 -1233 -549 -1229
rect -545 -1233 -536 -1229
rect -532 -1233 -526 -1229
rect -522 -1233 -516 -1229
rect -512 -1233 -504 -1229
rect -500 -1233 -492 -1229
rect -473 -1255 -468 -1206
rect -430 -1207 -306 -1204
rect -447 -1218 -421 -1213
rect -440 -1224 -436 -1218
rect -338 -1228 -334 -1207
rect -318 -1208 -306 -1207
rect -306 -1215 -294 -1211
rect -287 -1219 -279 -1197
rect -250 -1204 -246 -1141
rect -272 -1208 -246 -1204
rect -234 -1208 -230 -1047
rect -260 -1215 -240 -1211
rect -232 -1215 -230 -1208
rect -77 -1195 -71 -1191
rect -67 -1195 -61 -1191
rect -57 -1195 -47 -1191
rect -81 -1199 -77 -1195
rect -287 -1224 -149 -1219
rect -338 -1232 -294 -1228
rect -432 -1255 -428 -1244
rect -326 -1239 -306 -1235
rect -473 -1259 -439 -1255
rect -432 -1259 -361 -1255
rect -473 -1294 -468 -1259
rect -432 -1264 -428 -1259
rect -440 -1280 -436 -1274
rect -440 -1284 -428 -1280
rect -326 -1294 -321 -1239
rect -287 -1242 -279 -1224
rect -260 -1232 -240 -1228
rect -272 -1239 -250 -1235
rect -307 -1266 -303 -1262
rect -263 -1266 -259 -1262
rect -307 -1267 -259 -1266
rect -303 -1271 -297 -1267
rect -293 -1271 -285 -1267
rect -281 -1271 -273 -1267
rect -269 -1271 -263 -1267
rect -473 -1298 -321 -1294
rect -253 -1305 -250 -1239
rect -193 -1277 -189 -1224
rect -154 -1256 -149 -1224
rect -51 -1206 -47 -1195
rect -51 -1210 -44 -1206
rect -40 -1210 -25 -1206
rect -51 -1211 -25 -1210
rect -44 -1217 -40 -1211
rect -61 -1248 -57 -1239
rect -36 -1248 -32 -1237
rect -120 -1253 -69 -1249
rect -61 -1252 -43 -1248
rect -36 -1252 -25 -1248
rect -61 -1256 -57 -1252
rect -154 -1260 -81 -1256
rect -73 -1259 -57 -1256
rect -36 -1257 -32 -1252
rect -73 -1263 -65 -1259
rect -193 -1281 -175 -1277
rect -81 -1278 -77 -1273
rect -61 -1278 -57 -1273
rect -44 -1273 -40 -1267
rect -44 -1277 -39 -1273
rect -35 -1277 -32 -1273
rect -44 -1278 -41 -1277
rect -81 -1279 -41 -1278
rect -77 -1283 -71 -1279
rect -67 -1283 -61 -1279
rect -57 -1283 -41 -1279
rect -350 -1314 -237 -1305
<< m2contact >>
rect -439 649 -432 656
rect -326 647 -321 653
rect -439 555 -432 562
rect -315 543 -308 551
rect -242 547 -234 554
rect -185 655 -179 661
rect -363 503 -352 510
rect -242 528 -234 534
rect -362 448 -352 457
rect -439 149 -432 156
rect -326 147 -321 153
rect -439 55 -432 62
rect -315 43 -308 51
rect -242 47 -234 54
rect -185 155 -179 161
rect -363 3 -352 10
rect -242 28 -234 34
rect -362 -52 -352 -43
rect -440 -298 -433 -291
rect -312 -300 -306 -294
rect -440 -392 -433 -385
rect -316 -404 -309 -396
rect -243 -400 -235 -393
rect -364 -444 -353 -437
rect -243 -419 -235 -413
rect -363 -499 -353 -490
rect -438 -759 -431 -752
rect -317 -761 -311 -755
rect -438 -853 -431 -846
rect -314 -865 -307 -857
rect -241 -861 -233 -854
rect -362 -905 -351 -898
rect -241 -880 -233 -874
rect -361 -960 -351 -951
rect -437 -1113 -430 -1106
rect -322 -1115 -316 -1109
rect -437 -1207 -430 -1200
rect -313 -1219 -306 -1211
rect -240 -1215 -232 -1208
rect -361 -1259 -350 -1252
rect -240 -1234 -232 -1228
rect -127 -1253 -120 -1248
rect -360 -1314 -350 -1305
<< metal2 >>
rect -326 732 -175 737
rect -439 562 -432 649
rect -326 653 -321 732
rect -363 540 -308 543
rect -363 510 -352 540
rect -242 534 -234 547
rect -362 457 -352 503
rect -352 448 -351 454
rect -185 398 -179 655
rect -326 232 -175 237
rect -439 62 -432 149
rect -326 153 -321 232
rect -363 40 -308 43
rect -363 10 -352 40
rect -242 34 -234 47
rect -362 -43 -352 3
rect -352 -52 -351 -46
rect -185 -212 -179 155
rect -312 -218 -175 -212
rect -440 -385 -433 -298
rect -312 -294 -306 -218
rect -364 -407 -309 -404
rect -364 -437 -353 -407
rect -243 -413 -235 -400
rect -363 -490 -353 -444
rect -353 -499 -352 -493
rect -317 -721 -175 -715
rect -438 -846 -431 -759
rect -317 -755 -311 -721
rect -362 -868 -307 -865
rect -362 -898 -351 -868
rect -241 -874 -233 -861
rect -361 -951 -351 -905
rect -351 -960 -350 -954
rect -220 -1109 -214 -986
rect -437 -1200 -430 -1113
rect -316 -1115 -214 -1109
rect -220 -1180 -214 -1115
rect -220 -1186 -121 -1180
rect -361 -1222 -306 -1219
rect -361 -1252 -350 -1222
rect -240 -1228 -232 -1215
rect -127 -1248 -121 -1186
rect -360 -1305 -350 -1259
rect -350 -1314 -349 -1308
<< labels >>
rlabel metal1 -610 62 -608 64 3 clk
rlabel metal1 -543 34 -541 36 1 gnd
rlabel metal1 -543 97 -541 99 5 vdd
rlabel metal1 -558 97 -556 99 5 vdd
rlabel metal1 -599 97 -597 99 5 vdd
rlabel metal1 -598 34 -596 36 1 gnd
rlabel metal1 -499 34 -497 36 1 gnd
rlabel metal1 -499 97 -497 99 5 vdd
rlabel metal1 -610 55 -608 57 1 b3d
rlabel metal1 -491 61 -489 63 7 b3
rlabel metal1 -438 191 -433 192 1 gnd
rlabel metal1 -449 44 -423 49 5 vdd
rlabel metal1 -439 -21 -434 -20 1 gnd
rlabel metal1 -423 216 -421 218 7 a3bar
rlabel metal1 -425 4 -423 6 7 b3bar
rlabel metal1 -356 188 -330 193 5 vdd
rlabel metal1 -346 123 -341 124 1 gnd
rlabel metal1 -334 148 -332 150 7 g3
rlabel metal1 -281 111 -278 113 5 vdd
rlabel metal1 -281 -8 -278 -6 1 gnd
rlabel metal1 -217 39 -214 42 7 p3
rlabel metal1 -610 -283 -608 -281 3 clk
rlabel metal1 -543 -311 -541 -309 1 gnd
rlabel metal1 -543 -248 -541 -246 5 vdd
rlabel metal1 -558 -248 -556 -246 5 vdd
rlabel metal1 -599 -248 -597 -246 5 vdd
rlabel metal1 -598 -311 -596 -309 1 gnd
rlabel metal1 -499 -311 -497 -309 1 gnd
rlabel metal1 -499 -248 -497 -246 5 vdd
rlabel metal1 -610 -290 -608 -288 1 a2d
rlabel metal1 -491 -284 -489 -282 7 a2
rlabel metal1 -449 -191 -423 -186 5 vdd
rlabel metal1 -439 -256 -434 -255 1 gnd
rlabel metal1 -450 -403 -424 -398 5 vdd
rlabel metal1 -440 -468 -435 -467 1 gnd
rlabel metal1 -376 -261 -374 -260 1 vdd
rlabel metal1 -357 -259 -331 -254 5 vdd
rlabel metal1 -347 -324 -342 -323 1 gnd
rlabel metal1 -282 -336 -279 -334 5 vdd
rlabel metal1 -282 -455 -279 -453 1 gnd
rlabel metal1 -218 -408 -215 -405 7 p2
rlabel metal1 -335 -299 -332 -296 1 g2
rlabel metal1 -425 -232 -422 -229 1 a2bar
rlabel metal1 -426 -443 -423 -440 1 b2bar
rlabel metal1 -447 -652 -421 -647 5 vdd
rlabel metal1 -437 -717 -432 -716 1 gnd
rlabel metal1 -448 -864 -422 -859 5 vdd
rlabel metal1 -438 -929 -433 -928 1 gnd
rlabel metal1 -374 -722 -372 -721 1 vdd
rlabel metal1 -355 -720 -329 -715 5 vdd
rlabel metal1 -345 -785 -340 -784 1 gnd
rlabel metal1 -280 -797 -277 -795 5 vdd
rlabel metal1 -280 -916 -277 -914 1 gnd
rlabel metal1 -218 -869 -216 -867 7 p1
rlabel metal1 -333 -761 -329 -757 1 g1
rlabel metal1 -423 -693 -420 -690 1 a1bar
rlabel metal1 -424 -904 -421 -901 1 b1bar
rlabel metal1 -610 -847 -608 -845 3 clk
rlabel metal1 -543 -875 -541 -873 1 gnd
rlabel metal1 -543 -812 -541 -810 5 vdd
rlabel metal1 -558 -812 -556 -810 5 vdd
rlabel metal1 -599 -812 -597 -810 5 vdd
rlabel metal1 -598 -875 -596 -873 1 gnd
rlabel metal1 -499 -875 -497 -873 1 gnd
rlabel metal1 -499 -812 -497 -810 5 vdd
rlabel metal1 -610 -854 -608 -852 1 b1d
rlabel metal1 -491 -848 -489 -846 7 b1
rlabel metal1 -612 -744 -610 -742 3 clk
rlabel metal1 -545 -772 -543 -770 1 gnd
rlabel metal1 -545 -709 -543 -707 5 vdd
rlabel metal1 -560 -709 -558 -707 5 vdd
rlabel metal1 -601 -709 -599 -707 5 vdd
rlabel metal1 -600 -772 -598 -770 1 gnd
rlabel metal1 -501 -772 -499 -770 1 gnd
rlabel metal1 -501 -709 -499 -707 5 vdd
rlabel metal1 -493 -745 -491 -743 1 a1
rlabel metal1 -612 -751 -610 -749 1 a1d
rlabel metal1 -611 -385 -609 -383 3 clk
rlabel metal1 -544 -413 -542 -411 1 gnd
rlabel metal1 -544 -350 -542 -348 5 vdd
rlabel metal1 -559 -350 -557 -348 5 vdd
rlabel metal1 -600 -350 -598 -348 5 vdd
rlabel metal1 -599 -413 -597 -411 1 gnd
rlabel metal1 -500 -413 -498 -411 1 gnd
rlabel metal1 -500 -350 -498 -348 5 vdd
rlabel metal1 -611 -392 -609 -390 1 b2d
rlabel metal1 -492 -386 -490 -384 1 b2
rlabel metal1 -610 -1101 -608 -1099 3 a0d
rlabel metal1 -423 -1259 -419 -1255 1 b0bar
rlabel metal1 -422 -1047 -418 -1043 1 a0bar
rlabel metal1 -332 -1115 -328 -1111 1 g0
rlabel metal1 -279 -1151 -276 -1149 5 vdd
rlabel metal1 -344 -1139 -339 -1138 1 gnd
rlabel metal1 -354 -1074 -328 -1069 5 vdd
rlabel metal1 -373 -1076 -371 -1075 1 vdd
rlabel metal1 -437 -1283 -432 -1282 1 gnd
rlabel metal1 -447 -1218 -421 -1213 5 vdd
rlabel metal1 -436 -1071 -431 -1070 1 gnd
rlabel metal1 -446 -1006 -420 -1001 5 vdd
rlabel metal1 -609 -1211 -607 -1209 1 b0d
rlabel metal1 -490 -1205 -488 -1203 7 b0
rlabel metal1 -491 -1095 -489 -1093 7 a0
rlabel metal1 -498 -1169 -496 -1167 5 vdd
rlabel metal1 -498 -1232 -496 -1230 1 gnd
rlabel metal1 -597 -1232 -595 -1230 1 gnd
rlabel metal1 -598 -1169 -596 -1167 5 vdd
rlabel metal1 -557 -1169 -555 -1167 5 vdd
rlabel metal1 -542 -1169 -540 -1167 5 vdd
rlabel metal1 -542 -1232 -540 -1230 1 gnd
rlabel metal1 -609 -1204 -607 -1202 3 clk
rlabel metal1 -499 -1059 -497 -1057 5 vdd
rlabel metal1 -499 -1122 -497 -1120 1 gnd
rlabel metal1 -598 -1122 -596 -1120 1 gnd
rlabel metal1 -599 -1059 -597 -1057 5 vdd
rlabel metal1 -558 -1059 -556 -1057 5 vdd
rlabel metal1 -543 -1059 -541 -1057 5 vdd
rlabel metal1 -543 -1122 -541 -1120 1 gnd
rlabel metal1 -610 -1094 -608 -1092 3 clk
rlabel metal1 -448 256 -422 261 5 vdd
rlabel metal1 -375 186 -373 187 1 vdd
rlabel metal1 -608 157 -606 159 1 a3d
rlabel metal1 -489 163 -487 165 7 a3
rlabel metal1 -497 199 -495 201 5 vdd
rlabel metal1 -497 136 -495 138 1 gnd
rlabel metal1 -596 136 -594 138 1 gnd
rlabel metal1 -597 199 -595 201 5 vdd
rlabel metal1 -556 199 -554 201 5 vdd
rlabel metal1 -541 199 -539 201 5 vdd
rlabel metal1 -541 136 -539 138 1 gnd
rlabel metal1 -608 164 -606 166 3 clk
rlabel metal1 -610 562 -608 564 3 clk
rlabel metal1 -543 534 -541 536 1 gnd
rlabel metal1 -543 597 -541 599 5 vdd
rlabel metal1 -558 597 -556 599 5 vdd
rlabel metal1 -599 597 -597 599 5 vdd
rlabel metal1 -598 534 -596 536 1 gnd
rlabel metal1 -499 534 -497 536 1 gnd
rlabel metal1 -499 597 -497 599 5 vdd
rlabel metal1 -438 691 -433 692 1 gnd
rlabel metal1 -449 544 -423 549 5 vdd
rlabel metal1 -439 479 -434 480 1 gnd
rlabel metal1 -356 688 -330 693 5 vdd
rlabel metal1 -346 623 -341 624 1 gnd
rlabel metal1 -281 611 -278 613 5 vdd
rlabel metal1 -281 492 -278 494 1 gnd
rlabel metal1 -448 756 -422 761 5 vdd
rlabel metal1 -375 686 -373 687 1 vdd
rlabel metal1 -497 699 -495 701 5 vdd
rlabel metal1 -497 636 -495 638 1 gnd
rlabel metal1 -596 636 -594 638 1 gnd
rlabel metal1 -597 699 -595 701 5 vdd
rlabel metal1 -556 699 -554 701 5 vdd
rlabel metal1 -541 699 -539 701 5 vdd
rlabel metal1 -541 636 -539 638 1 gnd
rlabel metal1 -608 664 -606 666 3 clk
rlabel metal1 -609 656 -604 660 1 a4d
rlabel metal1 -491 663 -486 665 1 a4
rlabel metal1 -423 716 -421 718 1 a4bar
rlabel metal1 -334 648 -332 650 1 g4
rlabel metal1 -491 561 -489 563 1 b4
rlabel metal1 -610 555 -608 557 1 b4d
rlabel metal1 -425 504 -423 506 1 b4bar
rlabel metal1 -217 539 -214 542 1 p4
rlabel metal1 -279 -1270 -276 -1268 1 gnd
rlabel metal1 -217 -1223 -214 -1220 7 p0
rlabel metal1 -59 -1251 -57 -1249 1 nout
rlabel metal1 -65 -1194 -63 -1192 1 vdd
rlabel metal1 -65 -1282 -63 -1280 1 gnd
rlabel metal1 -30 -1250 -25 -1249 7 out
rlabel metal1 -86 -1252 -84 -1250 3 b
rlabel metal1 -86 -1259 -84 -1257 3 a
<< end >>
