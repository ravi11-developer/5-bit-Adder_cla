=================================

.include TSMC_180nm.txt
.option scale=90n

VDD  VDD  0     1.8

* Input A bus: A1-A5 with pulse patterns
VA1  A1   0     pulse 0 1.8 0 0.1n 0.1n 10n 20n
VA2  A2   0     pulse 0 1.8 0 0.1n 0.1n 20n 40n
VA3  A3   0     pulse 0 1.8 0 0.1n 0.1n 40n 80n
VA4  A4   0     pulse 0 1.8 0 0.1n 0.1n 80n 160n
VA5  A5   0     pulse 0 1.8 0 0.1n 0.1n 160n 320n

* Input B bus: B1-B5 with pulse patterns
VB1  B1   0     pulse 0 1.8 0 0.1n 0.1n 5n 10n
VB2  B2   0     pulse 0 1.8 0 0.1n 0.1n 15n 30n
VB3  B3   0     pulse 0 1.8 0 0.1n 0.1n 35n 70n
VB4  B4   0     pulse 0 1.8 0 0.1n 0.1n 75n 150n
VB5  B5   0     pulse 0 1.8 0 0.1n 0.1n 155n 310n

* Carry input
V_Cin  Cin  0 0

M1000 C2 P3 S3 w_663_115# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1001 C1 P2 S2 w_663_200# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1002 P4 B4 A4 w_2_72# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1003 C2 P2 C1 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1004 C3 P4 S4 w_672_28# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1005 C5 D5 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1006 a_671_213# P2 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1007 G1b A1 a_162_375# Gnd CMOSN w=8 l=2
+  ad=40p pd=26u as=24p ps=14u
M1008 Cin a_671_288# S1 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1009 a_278_n136# B1 D1 w_265_n142# CMOSP w=16 l=2
+  ad=48p pd=22u as=80p ps=42u
M1010 a_10_13# A5 VDD w_2_0# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1011 VDD A4 G4b w_281_395# CMOSP w=8 l=2
+  ad=40p pd=26u as=24p ps=14u
M1012 a_428_n136# B4 D4 w_415_n142# CMOSP w=16 l=2
+  ad=48p pd=22u as=80p ps=42u
M1013 G2b B2 VDD w_193_395# CMOSP w=8 l=2
+  ad=24p pd=14u as=40p ps=26u
M1014 C4 P5 S5 w_672_n108# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1015 C2 D2 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1016 C5 G5b VDD w_571_176# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1017 G1b B1 VDD w_149_395# CMOSP w=8 l=2
+  ad=24p pd=14u as=40p ps=26u
M1018 a_10_155# A3 VDD w_2_142# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1019 C3 P3b C2 w_362_176# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1020 P2 B2 A2 w_2_209# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1021 VDD A3 G3b w_237_395# CMOSP w=8 l=2
+  ad=40p pd=26u as=24p ps=14u
M1022 P1b P1 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1023 P5b P5 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1024 C5 P5 C4 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1025 B5 A5 P5 w_2_0# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1026 P3b P3 VDD w_54_186# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1027 C2 G2b VDD w_328_176# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1028 P5b P5 VDD w_54_44# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1029 a_680_n95# P5 VDD w_672_n108# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1030 S5 C4 a_680_n95# Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1031 a_10_13# A5 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1032 G5b A5 a_338_375# Gnd CMOSN w=8 l=2
+  ad=40p pd=26u as=24p ps=14u
M1033 a_250_375# B3 GND Gnd CMOSN w=8 l=2
+  ad=24p pd=14u as=40p ps=26u
M1034 P1 B1 A1 w_3_277# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1035 B3 A3 P3 w_2_142# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1036 VDD A1 a_278_n136# w_265_n142# CMOSP w=16 l=2
+  ad=80p pd=42u as=48p ps=22u
M1037 D1 B1 GND Gnd CMOSN w=4 l=2
+  ad=12p pd=10u as=20p ps=18u
M1038 S3 C2 P3 w_663_115# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1039 S2 C1 P2 w_663_200# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1040 VDD A4 a_428_n136# w_415_n142# CMOSP w=16 l=2
+  ad=80p pd=42u as=48p ps=22u
M1041 D4 B4 GND Gnd CMOSN w=4 l=2
+  ad=12p pd=10u as=20p ps=18u
M1042 C3 a_680_41# S4 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1043 a_380_n136# B3 D3 w_367_n142# CMOSP w=16 l=2
+  ad=48p pd=22u as=80p ps=42u
M1044 S4 C3 P4 w_672_28# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1045 P3 B3 a_10_155# Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1046 a_10_155# A3 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1047 B2 a_10_222# P2 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1048 P4b P4 VDD w_54_116# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1049 S1 Cin a_671_288# Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1050 G5b B5 VDD w_325_395# CMOSP w=8 l=2
+  ad=24p pd=14u as=40p ps=26u
M1051 C3 P3 C2 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1052 B4 A4 P4 w_2_72# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1053 a_671_288# P1 VDD w_663_275# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1054 G4b B4 VDD w_281_395# CMOSP w=8 l=2
+  ad=24p pd=14u as=40p ps=26u
M1055 B1 a_11_290# P1 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1056 P3b P3 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1057 C2 a_671_128# S3 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1058 C1 a_671_213# S2 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1059 P4 B4 a_10_85# Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1060 VDD A2 G2b w_193_395# CMOSP w=8 l=2
+  ad=40p pd=26u as=24p ps=14u
M1061 P5 B5 A5 w_2_0# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1062 P2b P2 VDD w_54_253# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1063 GND A1 D1 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=12p ps=10u
M1064 C3 D3 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1065 GND A4 D4 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=12p ps=10u
M1066 VDD A2 a_332_n136# w_319_n142# CMOSP w=16 l=2
+  ad=80p pd=42u as=48p ps=22u
M1067 S5 C4 P5 w_672_n108# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1068 B5 a_10_13# P5 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1069 VDD A3 a_380_n136# w_367_n142# CMOSP w=16 l=2
+  ad=80p pd=42u as=48p ps=22u
M1070 D3 B3 GND Gnd CMOSN w=4 l=2
+  ad=12p pd=10u as=20p ps=18u
M1071 a_487_n136# B5 D5 w_474_n142# CMOSP w=16 l=2
+  ad=48p pd=22u as=80p ps=42u
M1072 C4 P4b C3 w_443_176# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1073 VDD A1 G1b w_149_395# CMOSP w=8 l=2
+  ad=40p pd=26u as=24p ps=14u
M1074 G4b A4 a_294_375# Gnd CMOSN w=8 l=2
+  ad=40p pd=26u as=24p ps=14u
M1075 a_332_n136# B2 D2 w_319_n142# CMOSP w=16 l=2
+  ad=48p pd=22u as=80p ps=42u
M1076 a_671_128# P3 VDD w_663_115# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1077 a_206_375# B2 GND Gnd CMOSN w=8 l=2
+  ad=24p pd=14u as=40p ps=26u
M1078 P4b P4 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1079 C3 G3b VDD w_409_176# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1080 Cin P1 S1 w_663_275# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1081 a_671_288# P1 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1082 a_680_41# P4 VDD w_672_28# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1083 S4 C3 a_680_41# Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1084 a_10_85# A4 VDD w_2_72# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1085 P2 B2 a_10_222# Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1086 C1 P1b Cin w_200_176# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1087 a_162_375# B1 GND Gnd CMOSN w=8 l=2
+  ad=24p pd=14u as=40p ps=26u
M1088 G3b A3 a_250_375# Gnd CMOSN w=8 l=2
+  ad=40p pd=26u as=24p ps=14u
M1089 a_680_n95# P5 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1090 P1 B1 a_11_290# Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1091 GND A2 D2 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=12p ps=10u
M1092 B3 a_10_155# P3 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1093 P2b P2 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1094 GND A3 D3 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=12p ps=10u
M1095 S3 C2 a_671_128# Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1096 a_10_222# A2 VDD w_2_209# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1097 S2 C1 a_671_213# Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1098 VDD A5 a_487_n136# w_474_n142# CMOSP w=16 l=2
+  ad=80p pd=42u as=48p ps=22u
M1099 a_680_41# P4 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1100 a_671_128# P3 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1101 D5 B5 GND Gnd CMOSN w=4 l=2
+  ad=12p pd=10u as=20p ps=18u
M1102 C1 D1 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1103 C2 P2b C1 w_281_176# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1104 VDD A5 G5b w_325_395# CMOSP w=8 l=2
+  ad=40p pd=26u as=24p ps=14u
M1105 D2 B2 GND Gnd CMOSN w=4 l=2
+  ad=12p pd=10u as=20p ps=18u
M1106 G3b B3 VDD w_237_395# CMOSP w=8 l=2
+  ad=24p pd=14u as=40p ps=26u
M1107 a_10_85# A4 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1108 C4 P4 C3 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1109 a_11_290# A1 VDD w_3_277# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1110 P5 B5 a_10_13# Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1111 C4 a_680_n95# S5 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1112 C1 G1b VDD w_247_176# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1113 P3 B3 A3 w_2_142# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1114 B2 A2 P2 w_2_209# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1115 a_338_375# B5 GND Gnd CMOSN w=8 l=2
+  ad=24p pd=14u as=40p ps=26u
M1116 B4 a_10_85# P4 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1117 C1 P1 Cin Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1118 a_671_213# P2 VDD w_663_200# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1119 S1 Cin P1 w_663_275# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1120 C4 D4 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1121 P1b P1 VDD w_59_317# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1122 a_10_222# A2 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1123 a_294_375# B4 GND Gnd CMOSN w=8 l=2
+  ad=24p pd=14u as=40p ps=26u
M1124 C5 P5b C4 w_524_176# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1125 G2b A2 a_206_375# Gnd CMOSN w=8 l=2
+  ad=40p pd=26u as=24p ps=14u
M1126 B1 A1 P1 w_3_277# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1127 a_11_290# A1 GND Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1128 GND A5 D5 Gnd CMOSN w=4 l=2
+  ad=20p pd=18u as=12p ps=10u
M1129 C4 G4b VDD w_490_176# CMOSP w=8 l=2
+  ad=40p pd=26u as=40p ps=26u

C0 a_11_290# w_3_277# 0.00788f
C1 A4 P4 0.13929f
C2 a_487_n136# VDD 0.16495f
C3 w_524_176# C4 0.02413f
C4 a_10_222# B2 0.06848f
C5 w_281_176# G1b 0
C6 a_338_375# G5b 0.12374f
C7 P3 S3 0.13929f
C8 A4 VDD 0.10851f
C9 w_409_176# C3 0.00961f
C10 a_11_290# B1 0.06848f
C11 w_193_395# VDD 0.01594f
C12 w_281_395# B4 0.02415f
C13 C5 G5b 0.05805f
C14 D5 w_474_n142# 0.0095f
C15 G3b A3 0.01233f
C16 P4b D2 0.00115f
C17 G1b G3b 0.03324f
C18 P5b D1 0.00423f
C19 P1b VDD 0.08248f
C20 P2 GND 0.05686f
C21 D1 B1 0.00929f
C22 a_10_85# P4 0.16971f
C23 D1 w_265_n142# 0.0095f
C24 w_319_n142# A2 0.0261f
C25 w_663_200# VDD 0.01041f
C26 a_338_375# GND 0.08248f
C27 w_149_395# B1 0.02415f
C28 D2 P4 0.01433f
C29 P5b P5 0.11264f
C30 a_10_85# VDD 0.08248f
C31 a_680_n95# C4 0.06848f
C32 w_672_n108# a_680_n95# 0.00788f
C33 D4 a_428_n136# 0.16495f
C34 P1b P3b 0.01027f
C35 VDD A3 0.10851f
C36 G1b VDD 0.37467f
C37 a_206_375# GND 0.08248f
C38 C5 GND 0.0825f
C39 D4 B4 0.00929f
C40 P1b P1 0.09638f
C41 w_663_115# C2 0.04001f
C42 GND A2 0.00226f
C43 VDD a_680_n95# 0.08248f
C44 G2b A4 0
C45 w_474_n142# A5 0.0261f
C46 w_237_395# A3 0.02415f
C47 w_193_395# G2b 0.00809f
C48 w_200_176# P1b 0.05386f
C49 w_281_176# C2 0.00924f
C50 A5 P5 0.13929f
C51 GND a_10_13# 0.09279f
C52 a_10_155# B3 0.06848f
C53 P3b G1b 0.00876f
C54 w_490_176# P4b 0.00104f
C55 C1 P2b 0.18385f
C56 B4 P4 0.30607f
C57 a_428_n136# VDD 0.16495f
C58 w_490_176# C4 0.00961f
C59 w_247_176# G1b 0.05395f
C60 P3 a_671_128# 0.11618f
C61 B4 VDD 0.04965f
C62 w_2_142# A3 0.08314f
C63 w_362_176# C3 0.00924f
C64 Cin w_663_275# 0.04001f
C65 C5 D5 0.0566f
C66 a_671_213# VDD 0.08248f
C67 D3 A3 0.00182f
C68 w_490_176# VDD 0.01489f
C69 D2 G2b 0.00755f
C70 G2b A3 0
C71 G3b B3 0.00359f
C72 G1b G2b 0.06294f
C73 P5b C5 0.06743f
C74 Cin C1 0.29898f
C75 P4b D1 0
C76 a_10_222# GND 0.09279f
C77 D4 P5 0.01221f
C78 P3 C3 0.04196f
C79 a_11_290# VDD 0.08248f
C80 w_319_n142# B2 0.0261f
C81 w_54_253# VDD 0.00789f
C82 D1 P4 0.01221f
C83 a_294_375# GND 0.08248f
C84 C2 VDD 0.08248f
C85 a_680_n95# S5 0.11734f
C86 P5 C4 0.24159f
C87 w_672_n108# P5 0.08314f
C88 a_671_128# GND 0.09279f
C89 a_10_85# A4 0.11618f
C90 S4 C3 0.30607f
C91 VDD B3 0.04965f
C92 w_474_n142# VDD 0.00787f
C93 a_162_375# GND 0.08248f
C94 w_149_395# VDD 0.01594f
C95 C1 GND 0.0825f
C96 S2 w_663_200# 0.02113f
C97 a_11_290# P1 0.16405f
C98 w_663_115# S3 0.02113f
C99 C2 P3b 0.22478f
C100 GND B2 0.0025f
C101 VDD P5 0.05789f
C102 G2b B4 0
C103 w_474_n142# B5 0.0261f
C104 w_237_395# B3 0.02415f
C105 S1 w_663_275# 0.02113f
C106 A5 a_10_13# 0.11618f
C107 B5 P5 0.30607f
C108 GND C3 0.0825f
C109 w_443_176# G3b 0
C110 w_443_176# P4b 0.05377f
C111 P4b P2 0.00714f
C112 a_380_n136# VDD 0.16495f
C113 w_443_176# C4 0.00924f
C114 a_294_375# G4b 0.12374f
C115 w_2_142# B3 0.04001f
C116 C2 G2b 0.05905f
C117 B4 A4 0.49715f
C118 w_2_0# A5 0.08314f
C119 P2 VDD 0.05789f
C120 D3 B3 0.00929f
C121 D4 w_415_n142# 0.0095f
C122 G2b B3 0
C123 D3 P5 0.01221f
C124 P2b GND 0.09279f
C125 C5 C4 0.29898f
C126 w_2_209# VDD 0.01041f
C127 a_250_375# GND 0.08248f
C128 P2 P3b 0.01027f
C129 a_671_213# S2 0.11734f
C130 P5 S5 0.13929f
C131 C5 VDD 0.08248f
C132 D3 a_380_n136# 0.16495f
C133 a_10_85# B4 0.06848f
C134 P3 GND 0.05671f
C135 P1 P2 0.09247f
C136 a_680_41# C3 0.06848f
C137 VDD A2 0.10851f
C138 w_54_44# P5 0.02088f
C139 w_415_n142# VDD 0.00787f
C140 a_671_213# w_663_200# 0.00788f
C141 w_663_115# a_671_128# 0.00788f
C142 GND A1 0.00226f
C143 VDD a_10_13# 0.08248f
C144 a_671_288# w_663_275# 0.00788f
C145 w_571_176# C5 0.00961f
C146 B5 a_10_13# 0.06848f
C147 w_409_176# G3b 0.05395f
C148 w_281_176# C1 0.02413f
C149 Cin S1 0.30607f
C150 a_332_n136# VDD 0.16495f
C151 D2 C2 0.10666f
C152 w_2_0# VDD 0.01041f
C153 D5 G5b 0.00755f
C154 G2b a_206_375# 0.12374f
C155 w_3_277# A1 0.08314f
C156 w_409_176# VDD 0.01489f
C157 w_2_0# B5 0.04001f
C158 a_10_222# VDD 0.08248f
C159 D1 G1b 0.00755f
C160 B3 A3 0.49715f
C161 G2b A2 0.01233f
C162 D2 P5 0.01433f
C163 w_149_395# G1b 0.00811f
C164 B1 A1 0.49715f
C165 w_265_n142# A1 0.0261f
C166 G3b C3 0.05897f
C167 w_663_275# VDD 0.01041f
C168 P4b C3 0.18354f
C169 a_671_128# VDD 0.08248f
C170 P2 S2 0.13929f
C171 P5 a_680_n95# 0.11618f
C172 C3 C4 0.29898f
C173 C1 VDD 0.08248f
C174 D5 GND 0.285f
C175 w_281_176# P2b 0.05383f
C176 P4 C3 0.13769f
C177 a_680_41# S4 0.11734f
C178 VDD B2 0.04965f
C179 w_367_n142# VDD 0.00787f
C180 G5b A5 0.01233f
C181 P5b GND 0.09353f
C182 P2 w_663_200# 0.08314f
C183 P3 a_10_155# 0.18281f
C184 w_663_115# P3 0.08314f
C185 VDD C3 0.08248f
C186 GND B1 0.0025f
C187 w_415_n142# A4 0.0261f
C188 w_193_395# A2 0.02415f
C189 P1 w_663_275# 0.08314f
C190 w_524_176# C5 0.00924f
C191 w_54_116# P4b 0.00799f
C192 GND a_680_41# 0.09279f
C193 w_247_176# C1 0.00961f
C194 P3 w_54_186# 0.0209f
C195 C1 P1 0.04196f
C196 Cin a_671_288# 0.06848f
C197 a_278_n136# VDD 0.16495f
C198 w_54_116# P4 0.02088f
C199 P3b C3 0.05716f
C200 a_250_375# G3b 0.12374f
C201 w_200_176# C1 0.00924f
C202 A5 GND 0.00226f
C203 w_54_116# VDD 0.00789f
C204 G5b w_325_395# 0.00811f
C205 P4b P3 0.37646f
C206 w_3_277# B1 0.04001f
C207 a_10_155# GND 0.09279f
C208 D2 A2 0.00182f
C209 P2b VDD 0.08248f
C210 D3 w_367_n142# 0.0095f
C211 G2b B2 0.00359f
C212 D1 P5 0.01221f
C213 D3 C3 0.09229f
C214 a_671_288# GND 0.09279f
C215 w_265_n142# B1 0.0261f
C216 w_59_317# VDD 0.00789f
C217 P3 VDD 0.05789f
C218 P2b P3b 0.00876f
C219 P2 a_671_213# 0.11618f
C220 w_362_176# P3b 0.05383f
C221 w_672_28# C3 0.04001f
C222 G5b VDD 0.41507f
C223 D2 a_332_n136# 0.16495f
C224 D4 GND 0.28477f
C225 D5 A5 0.00182f
C226 a_671_288# S1 0.11734f
C227 P1 P2b 0.01027f
C228 P4 S4 0.13929f
C229 VDD A1 0.10851f
C230 G5b B5 0.00359f
C231 w_319_n142# VDD 0.00787f
C232 w_281_395# G4b 0.00811f
C233 P4b GND 0.09342f
C234 P2 w_54_253# 0.0209f
C235 C2 P2 0.04196f
C236 P3 P3b 0.09711f
C237 GND C4 0.0825f
C238 w_193_395# B2 0.02415f
C239 w_415_n142# B4 0.0261f
C240 w_571_176# G5b 0.05383f
C241 P1 w_59_317# 0.03264f
C242 D1 P2 0.01221f
C243 C1 S2 0.30607f
C244 GND P4 0.05744f
C245 w_362_176# G2b 0
C246 P3 w_2_142# 0.02113f
C247 C1 P1b 0.05716f
C248 Cin P1 0.24113f
C249 S3 C2 0.30607f
C250 w_2_72# P4 0.02113f
C251 P1 A1 0.13929f
C252 w_200_176# Cin 0.02413f
C253 C1 w_663_200# 0.04001f
C254 B5 GND 0.0025f
C255 w_2_72# VDD 0.01041f
C256 D4 G4b 0.00755f
C257 G1b a_162_375# 0.12374f
C258 P5b D4 0.00423f
C259 w_328_176# VDD 0.01489f
C260 D2 B2 0.00929f
C261 P3b GND 0.09279f
C262 C1 G1b 0.05897f
C263 G4b C4 0.05897f
C264 w_367_n142# A3 0.0261f
C265 P5b C4 0.18354f
C266 C5 P5 0.04196f
C267 P1 GND 0.02579f
C268 w_3_277# VDD 0.01041f
C269 a_10_13# P5 0.16971f
C270 w_672_28# S4 0.02113f
C271 G4b VDD 0.37467f
C272 w_325_395# A5 0.02415f
C273 P5b VDD 0.08248f
C274 D5 B5 0.00929f
C275 D3 GND 0.29513f
C276 P1 S1 0.13929f
C277 P1b P2b 0.01027f
C278 P4 a_680_41# 0.11618f
C279 VDD B1 0.04965f
C280 G2b GND 0
C281 w_265_n142# VDD 0.00787f
C282 P2 w_2_209# 0.02113f
C283 VDD a_680_41# 0.08248f
C284 P1b w_59_317# 0.00798f
C285 P1 w_3_277# 0.02113f
C286 C1 a_671_213# 0.06848f
C287 w_571_176# P5b 0.00157f
C288 w_2_0# P5 0.02113f
C289 P2 A2 0.13929f
C290 w_328_176# G2b 0.05398f
C291 P2b G1b 0.00876f
C292 Cin P1b 0.184f
C293 a_671_128# C2 0.06848f
C294 A5 VDD 0.10851f
C295 w_281_395# VDD 0.01594f
C296 P1 B1 0.30632f
C297 D2 P3 0.01433f
C298 C1 C2 0.29898f
C299 B5 A5 0.49715f
C300 A4 GND 0.00226f
C301 w_2_209# A2 0.08314f
C302 w_663_115# VDD 0.01041f
C303 a_10_155# VDD 0.08248f
C304 P3 A3 0.13929f
C305 P5b D3 0.00423f
C306 C1 D1 0.09218f
C307 G2b G4b 0.02475f
C308 w_2_72# A4 0.08314f
C309 C2 C3 0.29898f
C310 D4 C4 0.09828f
C311 a_671_288# VDD 0.08248f
C312 D2 w_319_n142# 0.0095f
C313 G1b A1 0.01233f
C314 w_367_n142# B3 0.0261f
C315 w_54_186# VDD 0.00789f
C316 P4b C4 0.06593f
C317 P1b GND 0.04124f
C318 w_672_n108# C4 0.04001f
C319 w_325_395# VDD 0.01594f
C320 P4b P4 0.18557f
C321 D5 a_487_n136# 0.16495f
C322 a_10_85# GND 0.09279f
C323 P5b w_54_44# 0.00802f
C324 a_10_222# P2 0.20331f
C325 P4 C4 0.04196f
C326 w_672_28# a_680_41# 0.00788f
C327 G3b VDD 0.37467f
C328 w_325_395# B5 0.02415f
C329 P4b VDD 0.08248f
C330 D1 a_278_n136# 0.16495f
C331 D2 GND 0.27446f
C332 P3b w_54_186# 0.00797f
C333 a_10_155# w_2_142# 0.00788f
C334 P1 a_671_288# 0.11618f
C335 w_2_72# a_10_85# 0.00788f
C336 VDD C4 0.08248f
C337 GND A3 0.00226f
C338 G2b A5 0
C339 G4b A4 0.01233f
C340 w_672_n108# VDD 0.01041f
C341 w_237_395# G3b 0.00811f
C342 P2b w_54_253# 0.00799f
C343 a_10_222# w_2_209# 0.00788f
C344 w_362_176# C2 0.02413f
C345 C2 P2b 0.05716f
C346 VDD P4 0.05789f
C347 GND a_680_n95# 0.09279f
C348 w_524_176# G4b 0
C349 w_524_176# P5b 0.05377f
C350 C1 P2 0.24125f
C351 P2 B2 0.30607f
C352 w_2_0# a_10_13# 0.00788f
C353 a_10_222# A2 0.11618f
C354 a_671_128# S3 0.11734f
C355 P3 C2 0.24154f
C356 B5 VDD 0.04965f
C357 a_11_290# A1 0.11618f
C358 w_443_176# C3 0.02413f
C359 w_237_395# VDD 0.01594f
C360 D1 P3 0.01221f
C361 D3 D4 0.05724f
C362 B4 GND 0.0025f
C363 w_2_209# B2 0.04001f
C364 w_571_176# VDD 0.01489f
C365 P3b VDD 0.08248f
C366 P3 B3 0.30607f
C367 w_281_395# A4 0.02415f
C368 D3 G3b 0.00755f
C369 P4b D3 0.00358f
C370 G2b G3b 0.02455f
C371 P5b D2 0.00498f
C372 a_671_213# GND 0.09279f
C373 D1 A1 0.00182f
C374 w_2_72# B4 0.04001f
C375 P1 VDD 0.09913f
C376 w_247_176# VDD 0.01489f
C377 B2 A2 0.49715f
C378 G1b B1 0.00359f
C379 w_149_395# A1 0.02415f
C380 a_11_290# GND 0.09279f
C381 D3 P4 0.01221f
C382 w_2_142# VDD 0.01041f
C383 S5 C4 0.30607f
C384 w_672_n108# S5 0.02113f
C385 C2 GND 0.0825f
C386 P1 P3b 0.01703f
C387 P2b P2 0.09711f
C388 w_672_28# P4 0.08314f
C389 G2b VDD 0.37483f
C390 D4 A4 0.00182f
C391 D1 GND 0.26415f
C392 GND B3 0.0025f
C393 w_672_28# VDD 0.01041f
C394 G2b B5 0
C395 G4b B4 0.00359f
C396 w_328_176# C2 0.00961f
C397 GND P5 0.05713f
C398 w_54_44# VDD 0.00789f
C399 a_10_155# A3 0.11618f
C400 w_490_176# G4b 0.05395f
C401 P3b G2b 0.01027f
C402 VDD 0 1.63268f
C403 a_487_n136# 0 0.00853f
C404 a_428_n136# 0 0.00853f
C405 a_380_n136# 0 0.00853f
C406 a_332_n136# 0 0.00853f
C407 a_278_n136# 0 0.00853f
C408 GND 0 1.39106f
C409 A5 0 0.71398f
C410 B5 0 0.53221f
C411 A4 0 0.71398f
C412 B4 0 0.53221f
C413 A3 0 0.71398f
C414 B3 0 0.53221f
C415 A2 0 0.71398f
C416 B2 0 0.53221f
C417 A1 0 0.71398f
C418 B1 0 0.53221f
C419 C4 0 0.69308f
C420 S5 0 0.3663f
C421 a_680_n95# 0 0.24503f
C422 P5 0 8.79655f
C423 a_10_13# 0 0.23914f
C424 C3 0 0.6764f
C425 S4 0 0.3663f
C426 a_680_41# 0 0.24503f
C427 P4 0 7.00365f
C428 a_10_85# 0 0.23914f
C429 C2 0 0.68616f
C430 S3 0 0.3663f
C431 a_671_128# 0 0.24503f
C432 P3 0 6.24858f
C433 D5 0 1.14244f
C434 D4 0 1.11908f
C435 D3 0 1.08724f
C436 D2 0 1.09833f
C437 D1 0 1.02853f
C438 C5 0 0.27082f
C439 C1 0 0.69015f
C440 Cin 0 0.45386f
C441 P5b 0 4.04682f
C442 P4b 0 2.54201f
C443 a_10_155# 0 0.23911f
C444 P3b 0 1.49444f
C445 S2 0 0.3663f
C446 a_671_213# 0 0.24503f
C447 P2 0 5.66891f
C448 a_10_222# 0 0.23909f
C449 P2b 0 1.72591f
C450 S1 0 0.3663f
C451 a_671_288# 0 0.24503f
C452 P1 0 5.66755f
C453 P1b 0 3.53543f
C454 a_11_290# 0 0.23919f
C455 a_338_375# 0 0.00433f
C456 a_294_375# 0 0.00433f
C457 a_250_375# 0 0.00433f
C458 a_206_375# 0 0.00433f
C459 a_162_375# 0 0.00433f
C460 G5b 0 1.80086f
C461 G4b 0 2.12344f
C462 G3b 0 2.33468f
C463 G2b 0 3.88162f
C464 G1b 0 2.62032f
C465 w_474_n142# 0 0.93208f
C466 w_415_n142# 0 0.93208f
C467 w_367_n142# 0 0.93208f
C468 w_319_n142# 0 0.93208f
C469 w_265_n142# 0 0.93208f
C470 w_672_n108# 0 1.25349f
C471 w_672_28# 0 1.25349f
C472 w_54_44# 0 0.48211f
C473 w_2_0# 0 1.25349f
C474 w_54_116# 0 0.48211f
C475 w_2_72# 0 1.25349f
C476 w_663_115# 0 1.25349f
C477 w_571_176# 0 0.67897f
C478 w_524_176# 0 0.67897f
C479 w_490_176# 0 0.67897f
C480 w_443_176# 0 0.67897f
C481 w_409_176# 0 0.67897f
C482 w_362_176# 0 0.67897f
C483 w_328_176# 0 0.67897f
C484 w_281_176# 0 0.67897f
C485 w_247_176# 0 0.67897f
C486 w_200_176# 0 0.67897f
C487 w_54_186# 0 0.48211f
C488 w_2_142# 0 1.25349f
C489 w_663_200# 0 1.25349f
C490 w_54_253# 0 0.48211f
C491 w_2_209# 0 1.25349f
C492 w_663_275# 0 1.25349f
C493 w_59_317# 0 0.48211f
C494 w_3_277# 0 1.25349f
C495 w_325_395# 0 0.64282f
C496 w_281_395# 0 0.64282f
C497 w_237_395# 0 0.64282f
C498 w_193_395# 0 0.64282f
C499 w_149_395# 0 0.64282f

.tran 0.01n 60n

* Propagation delay measurements
* Cin to S1 delay
.measure tran tpd_cin_s1_lh TRIG v(Cin) VAL=0.9 RISE=1 TARG v(S1) VAL=0.9 RISE=1
.measure tran tpd_cin_s1_hl TRIG v(Cin) VAL=0.9 FALL=1 TARG v(S1) VAL=0.9 FALL=1
.measure tran avg_tpd_cin_s1 param = '(tpd_cin_s1_lh + tpd_cin_s1_hl)/2'

* A1 to S1 delay
.measure tran tpd_a1_s1_lh TRIG v(A1) VAL=0.9 RISE=1 TARG v(S1) VAL=0.9 RISE=1
.measure tran tpd_a1_s1_hl TRIG v(A1) VAL=0.9 FALL=1 TARG v(S1) VAL=0.9 FALL=1
.measure tran avg_tpd_a1_s1 param = '(tpd_a1_s1_lh + tpd_a1_s1_hl)/2'

* B1 to S1 delay
.measure tran tpd_b1_s1_lh TRIG v(B1) VAL=0.9 RISE=1 TARG v(S1) VAL=0.9 RISE=1
.measure tran tpd_b1_s1_hl TRIG v(B1) VAL=0.9 FALL=1 TARG v(S1) VAL=0.9 FALL=1
.measure tran avg_tpd_b1_s1 param = '(tpd_b1_s1_lh + tpd_b1_s1_hl)/2'

* Cin to C1 delay (Carry propagation)
.measure tran tpd_cin_c1_lh TRIG v(Cin) VAL=0.9 RISE=1 TARG v(C1) VAL=0.9 RISE=1
.measure tran tpd_cin_c1_hl TRIG v(Cin) VAL=0.9 FALL=1 TARG v(C1) VAL=0.9 FALL=1
.measure tran avg_tpd_cin_c1 param = '(tpd_cin_c1_lh + tpd_cin_c1_hl)/2'

* A1 to C1 delay
.measure tran tpd_a1_c1_lh TRIG v(A1) VAL=0.9 RISE=1 TARG v(C1) VAL=0.9 RISE=1
.measure tran tpd_a1_c1_hl TRIG v(A1) VAL=0.9 FALL=1 TARG v(C1) VAL=0.9 FALL=1
.measure tran avg_tpd_a1_c1 param = '(tpd_a1_c1_lh + tpd_a1_c1_hl)/2'
.control
run
set hcopypscolor = 1
set color0=white
set xbrushwidth = 3
set curplottitle="2024102024_ravi__CLA_postlayout"

plot v(A1) v(B1)+2 v(C1)+4 v(S1)+6
plot v(A2) v(B2)+2 v(C2)+4 v(S2)+6
plot v(A3) v(B3)+2 v(C3)+4 v(S3)+6
plot v(A4) v(B4)+2 v(C4)+4 v(S4)+6
plot v(A5) v(B5)+2 v(C5)+4 v(S5)+6

* Print Sum outputs and Carry out
print v(S1) v(S2) v(S3) v(S4) v(S5) v(C5)

print delay_max
.endc
.end
