.include TSMC_180nm.txt
* Include TSMC 180nm technology file (model definitions for NMOS/PMOS)
.param SUPPLY=1.8
* Define supply voltage parameter = 1.8V
.option scale=90n
* Scale factor: all layout dimensions multiplied by 90nm
.global gnd vdd
* Global nodes: ground and power supply

Vdd vdd gnd 'SUPPLY'
* Voltage source: VDD = 1.8V
M1000 nout c vdd vdd CMOSP w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1001 a_n20_n101# e gnd Gnd CMOSN w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=0.11m
M1002 out nout gnd Gnd CMOSN w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1003 out nout vdd vdd CMOSP w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1004 nout e vdd vdd CMOSP w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1005 a_n8_n101# d a_n20_n101# Gnd CMOSN w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=60u
M1006 a_16_n101# b a_4_n101# Gnd CMOSN w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=60u
M1007 vdd b nout vdd CMOSP w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1008 a_4_n101# c a_n8_n101# Gnd CMOSN w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=60u
M1009 nout a a_16_n101# Gnd CMOSN w=50 l=2
+  ad=0.25n pd=0.11m as=0.25n ps=60u
M1010 nout a vdd vdd CMOSP w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1011 vdd d nout vdd CMOSP w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
C0 gnd a_16_n101# 1.13e-19
C1 gnd a_n20_n101# 1.13e-19
C2 a a_16_n101# 1.42e-19
C3 a a_n20_n101# 2.83e-19
C4 nout gnd 0.062834f
C5 c gnd 9.67e-19
C6 a nout 0.071424f
C7 c a 0.007761f
C8 d nout 0.083154f
C9 e b 0.007359f
C10 d c 0.341485f
C11 vdd a 0.020915f
C12 vdd d 0.020915f
C13 gnd a_n8_n101# 1.13e-19
C14 out gnd 0.130598f
C15 a a_n8_n101# 2.83e-19
C16 b gnd 9.67e-19
C17 e gnd 0.001936f
C18 b a 0.510277f
C19 c nout 0.008926f
C20 e a 0.007761f
C21 d b 0.007359f
C22 vdd nout 1.32495f
C23 vdd c 0.020915f
C24 e d 0.176533f
C25 gnd a_4_n101# 1.13e-19
C26 a a_4_n101# 2.83e-19
C27 a gnd 0.05598f
C28 nout out 0.060313f
C29 d gnd 9.67e-19
C30 b nout 0.008926f
C31 e nout 0.031122f
C32 c b 0.506518f
C33 d a 0.007761f
C34 vdd out 0.243018f
C35 vdd b 0.020915f
C36 e c 0.007278f
C37 vdd e 0.020698f
C38 gnd 0 0.736519f 
C39 out 0 0.105517f 
C40 nout 0 0.625451f 
C41 a 0 0.4646f 
C42 b 0 0.394239f 
C43 c 0 0.381196f 
C44 d 0 0.359481f 
C45 e 0 0.356293f 
C46 vdd 0 4.49066f 


va a gnd pulse 0 1.8 0 0.1n 0.1n 5n 10n
vb b gnd pulse 0 1.8 0 0.1n 0.1n 10n 20n
vc c gnd pulse 0 1.8 0 0.1n 0.1n 20n 40n
vd d gnd pulse 0 1.8 0 0.1n 0.1n 40n 80n
ve e gnd pulse 0 1.8 0 0.1n 0.1n 80n 160n

* Propagation delay measurements: inputs (a,b,c,d,e) -> out
.measure tran tpd_a_lh TRIG v(a) VAL=0.9 RISE=1 TARG v(out) VAL=0.9 RISE=1
.measure tran tpd_a_hl TRIG v(a) VAL=0.9 RISE=2 TARG v(out) VAL=0.9 FALL=1
.measure tran avg_tpd_a param = ((tpd_a_lh + tpd_a_hl)/2)

.measure tran tpd_b_lh TRIG v(b) VAL=0.9 RISE=1 TARG v(out) VAL=0.9 RISE=1
.measure tran tpd_b_hl TRIG v(b) VAL=0.9 RISE=2 TARG v(out) VAL=0.9 FALL=1
.measure tran avg_tpd_b param = ((tpd_b_lh + tpd_b_hl)/2)

.measure tran tpd_c_lh TRIG v(c) VAL=0.9 RISE=1 TARG v(out) VAL=0.9 RISE=1
.measure tran tpd_c_hl TRIG v(c) VAL=0.9 RISE=2 TARG v(out) VAL=0.9 FALL=1
.measure tran avg_tpd_c param = ((tpd_c_lh + tpd_c_hl)/2)

.measure tran tpd_d_lh TRIG v(d) VAL=0.9 RISE=1 TARG v(out) VAL=0.9 RISE=1
.measure tran tpd_d_hl TRIG v(d) VAL=0.9 RISE=2 TARG v(out) VAL=0.9 FALL=1
.measure tran avg_tpd_d param = ((tpd_d_lh + tpd_d_hl)/2)

.measure tran tpd_e_lh TRIG v(e) VAL=0.9 RISE=1 TARG v(out) VAL=0.9 RISE=1
.measure tran tpd_e_hl TRIG v(e) VAL=0.9 RISE=2 TARG v(out) VAL=0.9 FALL=1
.measure tran avg_tpd_e param = ((tpd_e_lh + tpd_e_hl)/2)

.tran 0.01n 200n

.control
run
set hcopypscolor = 1
set color0=white
set color1=black
plot v(a) v(b)+2 v(c)+4 v(d)+6 v(e)+8 v(out)+10
.endc