magic
tech scmos
timestamp 1763530775
<< nwell >>
rect -22 -29 26 48
<< ntransistor >>
rect -11 -69 -9 -59
rect 1 -69 3 -59
rect 13 -69 15 -59
<< ptransistor >>
rect -11 -23 -9 37
rect 1 -23 3 37
rect 13 -23 15 37
<< ndiffusion >>
rect -12 -69 -11 -59
rect -9 -69 -8 -59
rect 0 -69 1 -59
rect 3 -69 4 -59
rect 12 -69 13 -59
rect 15 -69 16 -59
<< pdiffusion >>
rect -12 -23 -11 37
rect -9 -23 1 37
rect 3 -23 13 37
rect 15 -23 16 37
<< ndcontact >>
rect -16 -69 -12 -59
rect -8 -69 0 -59
rect 4 -69 12 -59
rect 16 -69 20 -59
<< pdcontact >>
rect -16 -23 -12 37
rect 16 -23 20 37
<< psubstratepcontact >>
rect -16 -79 -12 -75
rect -6 -79 -2 -75
rect 6 -79 10 -75
rect 16 -79 20 -75
<< nsubstratencontact >>
rect -16 41 -12 45
rect -7 41 -3 45
rect 5 41 9 45
rect 16 41 20 45
<< polysilicon >>
rect -11 37 -9 40
rect 1 37 3 40
rect 13 37 15 40
rect -11 -59 -9 -23
rect 1 -59 3 -23
rect 13 -59 15 -23
rect -11 -72 -9 -69
rect 1 -72 3 -69
rect 13 -72 15 -69
<< polycontact >>
rect -16 -35 -11 -31
rect -4 -42 1 -38
rect 8 -49 13 -45
<< metal1 >>
rect -12 41 -7 45
rect -3 41 5 45
rect 9 41 16 45
rect 20 41 26 45
rect -16 37 -12 41
rect 16 -30 20 -23
rect -22 -35 -16 -31
rect 16 -34 26 -30
rect -22 -42 -4 -38
rect -22 -49 8 -45
rect 16 -52 20 -34
rect -8 -56 20 -52
rect -8 -59 0 -56
rect 16 -59 20 -56
rect -16 -74 -12 -69
rect 4 -74 12 -69
rect -16 -75 20 -74
rect -12 -79 -6 -75
rect -2 -79 6 -75
rect 10 -79 16 -75
<< labels >>
rlabel metal1 -22 -48 -20 -46 3 c
rlabel metal1 -21 -41 -19 -39 3 b
rlabel metal1 -21 -34 -19 -32 3 a
rlabel metal1 -1 42 2 44 5 vdd
rlabel metal1 17 -33 19 -31 1 nout
rlabel metal1 0 -78 2 -76 1 gnd
<< end >>
