magic
tech scmos
timestamp 1764769537
<< nwell >>
rect -20 84 86 183
rect -20 65 98 84
rect 72 44 98 65
<< ntransistor >>
rect 84 21 86 31
rect -8 9 -5 19
rect 11 9 13 19
rect 23 9 25 19
rect 35 9 37 19
rect 47 9 49 19
rect 59 9 61 19
<< ptransistor >>
rect -8 71 -5 171
rect 11 71 13 171
rect 23 71 25 171
rect 35 71 37 171
rect 47 71 49 171
rect 59 71 61 171
rect 84 51 86 71
<< ndiffusion >>
rect 83 21 84 31
rect 86 21 87 31
rect -9 9 -8 19
rect -5 9 -3 19
rect 10 9 11 19
rect 13 9 14 19
rect 22 9 23 19
rect 25 9 26 19
rect 34 9 35 19
rect 37 9 38 19
rect 46 9 47 19
rect 49 9 50 19
rect 58 9 59 19
rect 61 9 62 19
<< pdiffusion >>
rect -9 71 -8 171
rect -5 71 11 171
rect 13 71 23 171
rect 25 71 35 171
rect 37 71 47 171
rect 49 71 59 171
rect 61 71 62 171
rect 83 51 84 71
rect 86 51 87 71
<< ndcontact >>
rect 79 21 83 31
rect 87 21 91 31
rect -13 9 -9 19
rect -3 9 10 19
rect 14 9 22 19
rect 26 9 34 19
rect 38 9 46 19
rect 50 9 58 19
rect 62 9 66 19
<< pdcontact >>
rect -13 71 -9 171
rect 62 71 66 171
rect 79 51 83 71
rect 87 51 91 71
<< psubstratepcontact >>
rect -1 1 4 5
rect 16 0 20 4
rect 27 1 31 5
rect 40 0 44 4
rect 52 0 56 4
rect 79 8 83 12
rect 62 0 66 4
<< nsubstratencontact >>
rect 4 176 10 180
rect 15 176 21 180
rect 27 176 32 180
rect 39 176 45 180
rect 52 176 58 180
rect 63 176 67 180
rect 79 83 83 87
<< polysilicon >>
rect -8 171 -5 186
rect 11 171 13 186
rect 23 171 25 186
rect 35 171 37 186
rect 47 171 49 186
rect 59 171 61 186
rect 84 71 86 74
rect -8 19 -5 71
rect 11 19 13 71
rect 23 19 25 71
rect 35 19 37 71
rect 47 19 49 71
rect 59 19 61 71
rect 84 31 86 51
rect 84 16 86 21
rect -8 -2 -5 9
rect 11 -2 13 9
rect 23 -2 25 9
rect 35 -2 37 9
rect 47 -2 49 9
rect 59 -2 61 9
<< polycontact >>
rect -12 58 -8 62
rect 7 58 11 62
rect 19 51 23 55
rect 31 44 35 48
rect 43 37 47 41
rect 55 30 59 34
rect 80 36 84 40
<< metal1 >>
rect -13 180 83 181
rect -13 176 4 180
rect 10 176 15 180
rect 21 176 27 180
rect 32 176 39 180
rect 45 176 52 180
rect 58 176 63 180
rect 67 176 83 180
rect -13 175 83 176
rect -13 171 -9 175
rect -17 58 -12 62
rect 0 58 7 62
rect 0 51 19 55
rect 0 44 31 48
rect 0 37 43 41
rect 62 40 66 71
rect 79 87 83 175
rect 79 71 83 83
rect 87 40 91 51
rect 62 36 80 40
rect 87 36 98 40
rect 0 30 55 34
rect 62 27 66 36
rect 87 31 91 36
rect -13 22 66 27
rect -13 19 -9 22
rect 14 19 22 22
rect 38 19 46 22
rect 62 19 66 22
rect 79 12 83 21
rect -3 5 10 9
rect 26 5 34 9
rect 50 5 58 9
rect 79 5 83 8
rect -3 1 -1 5
rect 4 4 27 5
rect 4 1 16 4
rect -3 0 16 1
rect 20 1 27 4
rect 31 4 83 5
rect 31 1 40 4
rect 20 0 40 1
rect 44 0 52 4
rect 56 0 62 4
rect 66 0 83 4
<< labels >>
rlabel metal1 34 1 37 3 1 gnd
rlabel metal1 2 31 5 33 3 a
rlabel metal1 2 38 5 40 3 b
rlabel metal1 2 45 5 47 3 c
rlabel metal1 2 52 5 54 3 d
rlabel metal1 2 59 5 61 3 e
rlabel metal1 34 177 37 179 5 vdd
rlabel metal1 93 38 98 39 7 out
rlabel metal1 63 37 65 39 1 nout
rlabel metal1 -16 59 -14 61 3 f
<< end >>
