magic
tech scmos
timestamp 1764875535
<< nwell >>
rect 1328 944 1452 981
rect -448 623 -422 657
rect -609 568 -485 605
rect -392 555 -330 598
rect -145 579 -83 622
rect 365 586 471 712
rect 962 593 988 627
rect 365 567 483 586
rect 457 546 483 567
rect 1091 564 1151 622
rect 1322 558 1446 595
rect -611 466 -487 503
rect -315 459 -255 517
rect -72 485 -10 528
rect 964 477 990 511
rect -449 411 -423 445
rect 14 384 76 427
rect 119 364 181 407
rect 245 305 307 348
rect -448 223 -422 257
rect -609 168 -485 205
rect -392 155 -330 198
rect -112 172 -50 215
rect 357 174 443 273
rect 962 193 988 227
rect 357 155 455 174
rect 1091 164 1151 222
rect 1322 158 1446 195
rect 429 134 455 155
rect -611 66 -487 103
rect -315 59 -255 117
rect 7 91 69 134
rect 964 77 990 111
rect -449 11 -423 45
rect 122 -5 184 38
rect 250 -92 312 -49
rect -449 -224 -423 -190
rect -611 -279 -487 -242
rect -393 -292 -331 -249
rect -115 -273 -53 -230
rect 303 -289 389 -192
rect 953 -265 979 -231
rect 1082 -294 1142 -236
rect -612 -381 -488 -344
rect -316 -388 -256 -330
rect 16 -345 78 -302
rect 1319 -303 1443 -266
rect 955 -381 981 -347
rect -450 -436 -424 -402
rect 159 -428 221 -385
rect -447 -685 -421 -651
rect -613 -740 -489 -703
rect -391 -753 -329 -710
rect -94 -782 -32 -739
rect 127 -756 201 -682
rect 127 -759 175 -756
rect 915 -774 941 -740
rect -611 -843 -487 -806
rect -314 -849 -254 -791
rect 1044 -803 1104 -745
rect -448 -897 -422 -863
rect 7 -874 69 -831
rect 1322 -839 1446 -802
rect 917 -890 943 -856
rect -693 -1047 -569 -1010
rect -446 -1139 -420 -1105
rect -611 -1190 -487 -1153
rect -390 -1207 -328 -1164
rect -121 -1189 -59 -1146
rect 891 -1197 917 -1163
rect 1020 -1226 1080 -1168
rect -610 -1300 -486 -1263
rect -313 -1303 -253 -1245
rect -6 -1252 58 -1227
rect 1314 -1249 1438 -1212
rect -6 -1285 57 -1252
rect -6 -1286 31 -1285
rect 893 -1313 919 -1279
rect -447 -1351 -421 -1317
<< ntransistor >>
rect 1339 919 1341 929
rect 1374 919 1376 929
rect 1386 919 1388 929
rect 1407 919 1409 929
rect 1419 919 1421 929
rect 1439 919 1441 929
rect -436 600 -434 610
rect -598 543 -596 553
rect -563 543 -561 553
rect -551 543 -549 553
rect -530 543 -528 553
rect -518 543 -516 553
rect -498 543 -496 553
rect -381 516 -379 536
rect -369 516 -367 536
rect -344 532 -342 542
rect -134 540 -132 560
rect -122 540 -120 560
rect -97 556 -95 566
rect -600 441 -598 451
rect 974 570 976 580
rect 469 523 471 533
rect 1333 533 1335 543
rect 377 501 380 511
rect 396 501 398 511
rect 408 501 410 511
rect 420 501 422 511
rect 432 501 434 511
rect 444 501 446 511
rect 1102 505 1104 525
rect 1114 505 1116 525
rect 1126 505 1128 525
rect 1138 505 1140 525
rect 1368 533 1370 543
rect 1380 533 1382 543
rect 1401 533 1403 543
rect 1413 533 1415 543
rect 1433 533 1435 543
rect -565 441 -563 451
rect -553 441 -551 451
rect -532 441 -530 451
rect -520 441 -518 451
rect -500 441 -498 451
rect -61 446 -59 466
rect -49 446 -47 466
rect -24 462 -22 472
rect 976 454 978 464
rect -304 400 -302 420
rect -292 400 -290 420
rect -280 400 -278 420
rect -268 400 -266 420
rect -437 388 -435 398
rect 25 345 27 365
rect 37 345 39 365
rect 62 361 64 371
rect 130 325 132 345
rect 142 325 144 345
rect 167 341 169 351
rect 256 266 258 286
rect 268 266 270 286
rect 293 282 295 292
rect -436 200 -434 210
rect -598 143 -596 153
rect -563 143 -561 153
rect -551 143 -549 153
rect -530 143 -528 153
rect -518 143 -516 153
rect -498 143 -496 153
rect 974 170 976 180
rect -381 116 -379 136
rect -369 116 -367 136
rect -344 132 -342 142
rect -101 133 -99 153
rect -89 133 -87 153
rect -64 149 -62 159
rect -600 41 -598 51
rect 1333 133 1335 143
rect 441 111 443 121
rect 368 99 370 109
rect 380 99 382 109
rect 392 99 394 109
rect 404 99 406 109
rect 416 99 418 109
rect 1102 105 1104 125
rect 1114 105 1116 125
rect 1126 105 1128 125
rect 1138 105 1140 125
rect 1368 133 1370 143
rect 1380 133 1382 143
rect 1401 133 1403 143
rect 1413 133 1415 143
rect 1433 133 1435 143
rect -565 41 -563 51
rect -553 41 -551 51
rect -532 41 -530 51
rect -520 41 -518 51
rect -500 41 -498 51
rect 18 52 20 72
rect 30 52 32 72
rect 55 68 57 78
rect 976 54 978 64
rect -304 0 -302 20
rect -292 0 -290 20
rect -280 0 -278 20
rect -268 0 -266 20
rect -437 -12 -435 -2
rect 133 -44 135 -24
rect 145 -44 147 -24
rect 170 -28 172 -18
rect 261 -131 263 -111
rect 273 -131 275 -111
rect 298 -115 300 -105
rect -437 -247 -435 -237
rect -600 -304 -598 -294
rect -565 -304 -563 -294
rect -553 -304 -551 -294
rect -532 -304 -530 -294
rect -520 -304 -518 -294
rect -500 -304 -498 -294
rect -382 -331 -380 -311
rect -370 -331 -368 -311
rect -345 -315 -343 -305
rect -104 -312 -102 -292
rect -92 -312 -90 -292
rect -67 -296 -65 -286
rect 965 -288 967 -278
rect 375 -312 377 -302
rect 314 -332 316 -322
rect 326 -332 328 -322
rect 338 -332 340 -322
rect 350 -332 352 -322
rect 1330 -328 1332 -318
rect -601 -406 -599 -396
rect 1093 -353 1095 -333
rect 1105 -353 1107 -333
rect 1117 -353 1119 -333
rect 1129 -353 1131 -333
rect 1365 -328 1367 -318
rect 1377 -328 1379 -318
rect 1398 -328 1400 -318
rect 1410 -328 1412 -318
rect 1430 -328 1432 -318
rect -566 -406 -564 -396
rect -554 -406 -552 -396
rect -533 -406 -531 -396
rect -521 -406 -519 -396
rect -501 -406 -499 -396
rect 27 -384 29 -364
rect 39 -384 41 -364
rect 64 -368 66 -358
rect 967 -404 969 -394
rect -305 -447 -303 -427
rect -293 -447 -291 -427
rect -281 -447 -279 -427
rect -269 -447 -267 -427
rect -438 -459 -436 -449
rect 170 -467 172 -447
rect 182 -467 184 -447
rect 207 -451 209 -441
rect -435 -708 -433 -698
rect -602 -765 -600 -755
rect -567 -765 -565 -755
rect -555 -765 -553 -755
rect -534 -765 -532 -755
rect -522 -765 -520 -755
rect -502 -765 -500 -755
rect -380 -792 -378 -772
rect -368 -792 -366 -772
rect -343 -776 -341 -766
rect 187 -779 189 -769
rect -600 -868 -598 -858
rect -83 -821 -81 -801
rect -71 -821 -69 -801
rect -46 -805 -44 -795
rect 138 -799 140 -789
rect 150 -799 152 -789
rect 162 -799 164 -789
rect 927 -797 929 -787
rect -565 -868 -563 -858
rect -553 -868 -551 -858
rect -532 -868 -530 -858
rect -520 -868 -518 -858
rect -500 -868 -498 -858
rect 1055 -862 1057 -842
rect 1067 -862 1069 -842
rect 1079 -862 1081 -842
rect 1091 -862 1093 -842
rect -303 -908 -301 -888
rect -291 -908 -289 -888
rect -279 -908 -277 -888
rect -267 -908 -265 -888
rect 1333 -864 1335 -854
rect 1368 -864 1370 -854
rect 1380 -864 1382 -854
rect 1401 -864 1403 -854
rect 1413 -864 1415 -854
rect 1433 -864 1435 -854
rect -436 -920 -434 -910
rect 18 -913 20 -893
rect 30 -913 32 -893
rect 55 -897 57 -887
rect 929 -913 931 -903
rect -682 -1072 -680 -1062
rect -647 -1072 -645 -1062
rect -635 -1072 -633 -1062
rect -614 -1072 -612 -1062
rect -602 -1072 -600 -1062
rect -582 -1072 -580 -1062
rect -434 -1162 -432 -1152
rect -600 -1215 -598 -1205
rect -565 -1215 -563 -1205
rect -553 -1215 -551 -1205
rect -532 -1215 -530 -1205
rect -520 -1215 -518 -1205
rect -500 -1215 -498 -1205
rect -379 -1246 -377 -1226
rect -367 -1246 -365 -1226
rect -342 -1230 -340 -1220
rect -110 -1228 -108 -1208
rect -98 -1228 -96 -1208
rect -73 -1212 -71 -1202
rect 903 -1220 905 -1210
rect -599 -1325 -597 -1315
rect -564 -1325 -562 -1315
rect -552 -1325 -550 -1315
rect -531 -1325 -529 -1315
rect -519 -1325 -517 -1315
rect -499 -1325 -497 -1315
rect 1031 -1285 1033 -1265
rect 1043 -1285 1045 -1265
rect 1055 -1285 1057 -1265
rect 1067 -1285 1069 -1265
rect 1325 -1274 1327 -1264
rect 6 -1314 8 -1304
rect 18 -1314 20 -1304
rect 43 -1308 45 -1298
rect 1360 -1274 1362 -1264
rect 1372 -1274 1374 -1264
rect 1393 -1274 1395 -1264
rect 1405 -1274 1407 -1264
rect 1425 -1274 1427 -1264
rect 905 -1336 907 -1326
rect -302 -1362 -300 -1342
rect -290 -1362 -288 -1342
rect -278 -1362 -276 -1342
rect -266 -1362 -264 -1342
rect -435 -1374 -433 -1364
<< ptransistor >>
rect 1339 950 1341 970
rect 1351 950 1353 970
rect 1374 950 1376 970
rect 1407 950 1409 970
rect 1439 950 1441 970
rect -436 630 -434 650
rect -598 574 -596 594
rect -586 574 -584 594
rect -563 574 -561 594
rect -530 574 -528 594
rect -498 574 -496 594
rect -134 585 -132 605
rect -122 585 -120 605
rect -97 586 -95 606
rect -381 561 -379 581
rect -369 561 -367 581
rect -344 562 -342 582
rect 377 573 380 699
rect 396 573 398 699
rect 408 573 410 699
rect 420 573 422 699
rect 432 573 434 699
rect 444 573 446 699
rect 974 600 976 620
rect -600 472 -598 492
rect -588 472 -586 492
rect -565 472 -563 492
rect -532 472 -530 492
rect -500 472 -498 492
rect -304 465 -302 505
rect -292 465 -290 505
rect -280 465 -278 505
rect -268 465 -266 505
rect -61 491 -59 511
rect -49 491 -47 511
rect -24 492 -22 512
rect 469 553 471 573
rect 1102 570 1104 610
rect 1114 570 1116 610
rect 1126 570 1128 610
rect 1138 570 1140 610
rect 1333 564 1335 584
rect 1345 564 1347 584
rect 1368 564 1370 584
rect 1401 564 1403 584
rect 1433 564 1435 584
rect 976 484 978 504
rect -437 418 -435 438
rect 25 390 27 410
rect 37 390 39 410
rect 62 391 64 411
rect 130 370 132 390
rect 142 370 144 390
rect 167 371 169 391
rect 256 311 258 331
rect 268 311 270 331
rect 293 312 295 332
rect -436 230 -434 250
rect -598 174 -596 194
rect -586 174 -584 194
rect -563 174 -561 194
rect -530 174 -528 194
rect -498 174 -496 194
rect -381 161 -379 181
rect -369 161 -367 181
rect -344 162 -342 182
rect -101 178 -99 198
rect -89 178 -87 198
rect -64 179 -62 199
rect 368 161 370 261
rect 380 161 382 261
rect 392 161 394 261
rect 404 161 406 261
rect 416 161 418 261
rect 974 200 976 220
rect 1102 170 1104 210
rect 1114 170 1116 210
rect 1126 170 1128 210
rect 1138 170 1140 210
rect -600 72 -598 92
rect -588 72 -586 92
rect -565 72 -563 92
rect -532 72 -530 92
rect -500 72 -498 92
rect -304 65 -302 105
rect -292 65 -290 105
rect -280 65 -278 105
rect -268 65 -266 105
rect 18 97 20 117
rect 30 97 32 117
rect 55 98 57 118
rect 441 141 443 161
rect 1333 164 1335 184
rect 1345 164 1347 184
rect 1368 164 1370 184
rect 1401 164 1403 184
rect 1433 164 1435 184
rect 976 84 978 104
rect -437 18 -435 38
rect 133 1 135 21
rect 145 1 147 21
rect 170 2 172 22
rect 261 -86 263 -66
rect 273 -86 275 -66
rect 298 -85 300 -65
rect -437 -217 -435 -197
rect -600 -273 -598 -253
rect -588 -273 -586 -253
rect -565 -273 -563 -253
rect -532 -273 -530 -253
rect -500 -273 -498 -253
rect -382 -286 -380 -266
rect -370 -286 -368 -266
rect -345 -285 -343 -265
rect -104 -267 -102 -247
rect -92 -267 -90 -247
rect -67 -266 -65 -246
rect 314 -283 316 -203
rect 326 -283 328 -203
rect 338 -283 340 -203
rect 350 -283 352 -203
rect 965 -258 967 -238
rect 375 -282 377 -262
rect 27 -339 29 -319
rect 39 -339 41 -319
rect 64 -338 66 -318
rect 1093 -288 1095 -248
rect 1105 -288 1107 -248
rect 1117 -288 1119 -248
rect 1129 -288 1131 -248
rect 1330 -297 1332 -277
rect 1342 -297 1344 -277
rect 1365 -297 1367 -277
rect 1398 -297 1400 -277
rect 1430 -297 1432 -277
rect -601 -375 -599 -355
rect -589 -375 -587 -355
rect -566 -375 -564 -355
rect -533 -375 -531 -355
rect -501 -375 -499 -355
rect -305 -382 -303 -342
rect -293 -382 -291 -342
rect -281 -382 -279 -342
rect -269 -382 -267 -342
rect 967 -374 969 -354
rect -438 -429 -436 -409
rect 170 -422 172 -402
rect 182 -422 184 -402
rect 207 -421 209 -401
rect -435 -678 -433 -658
rect -602 -734 -600 -714
rect -590 -734 -588 -714
rect -567 -734 -565 -714
rect -534 -734 -532 -714
rect -502 -734 -500 -714
rect -380 -747 -378 -727
rect -368 -747 -366 -727
rect -343 -746 -341 -726
rect 138 -753 140 -693
rect 150 -753 152 -693
rect 162 -753 164 -693
rect 187 -749 189 -729
rect -83 -776 -81 -756
rect -71 -776 -69 -756
rect -46 -775 -44 -755
rect 927 -767 929 -747
rect -600 -837 -598 -817
rect -588 -837 -586 -817
rect -565 -837 -563 -817
rect -532 -837 -530 -817
rect -500 -837 -498 -817
rect -303 -843 -301 -803
rect -291 -843 -289 -803
rect -279 -843 -277 -803
rect -267 -843 -265 -803
rect 1055 -797 1057 -757
rect 1067 -797 1069 -757
rect 1079 -797 1081 -757
rect 1091 -797 1093 -757
rect 1333 -833 1335 -813
rect 1345 -833 1347 -813
rect 1368 -833 1370 -813
rect 1401 -833 1403 -813
rect 1433 -833 1435 -813
rect 18 -868 20 -848
rect 30 -868 32 -848
rect 55 -867 57 -847
rect -436 -890 -434 -870
rect 929 -883 931 -863
rect -682 -1041 -680 -1021
rect -670 -1041 -668 -1021
rect -647 -1041 -645 -1021
rect -614 -1041 -612 -1021
rect -582 -1041 -580 -1021
rect -434 -1132 -432 -1112
rect -600 -1184 -598 -1164
rect -588 -1184 -586 -1164
rect -565 -1184 -563 -1164
rect -532 -1184 -530 -1164
rect -500 -1184 -498 -1164
rect -379 -1201 -377 -1181
rect -367 -1201 -365 -1181
rect -342 -1200 -340 -1180
rect -110 -1183 -108 -1163
rect -98 -1183 -96 -1163
rect -73 -1182 -71 -1162
rect 903 -1190 905 -1170
rect 1031 -1220 1033 -1180
rect 1043 -1220 1045 -1180
rect 1055 -1220 1057 -1180
rect 1067 -1220 1069 -1180
rect -599 -1294 -597 -1274
rect -587 -1294 -585 -1274
rect -564 -1294 -562 -1274
rect -531 -1294 -529 -1274
rect -499 -1294 -497 -1274
rect -302 -1297 -300 -1257
rect -290 -1297 -288 -1257
rect -278 -1297 -276 -1257
rect -266 -1297 -264 -1257
rect 6 -1280 8 -1240
rect 18 -1280 20 -1240
rect 1325 -1243 1327 -1223
rect 1337 -1243 1339 -1223
rect 1360 -1243 1362 -1223
rect 1393 -1243 1395 -1223
rect 1425 -1243 1427 -1223
rect 43 -1278 45 -1258
rect 905 -1306 907 -1286
rect -435 -1344 -433 -1324
<< ndiffusion >>
rect 1338 919 1339 929
rect 1341 919 1342 929
rect 1373 919 1374 929
rect 1376 919 1386 929
rect 1388 919 1389 929
rect 1406 919 1407 929
rect 1409 919 1419 929
rect 1421 919 1422 929
rect 1438 919 1439 929
rect 1441 919 1442 929
rect -437 600 -436 610
rect -434 600 -433 610
rect -599 543 -598 553
rect -596 543 -595 553
rect -564 543 -563 553
rect -561 543 -551 553
rect -549 543 -548 553
rect -531 543 -530 553
rect -528 543 -518 553
rect -516 543 -515 553
rect -499 543 -498 553
rect -496 543 -495 553
rect -382 516 -381 536
rect -379 516 -369 536
rect -367 516 -366 536
rect -345 532 -344 542
rect -342 532 -341 542
rect -135 540 -134 560
rect -132 540 -122 560
rect -120 540 -119 560
rect -98 556 -97 566
rect -95 556 -94 566
rect -601 441 -600 451
rect -598 441 -597 451
rect 973 570 974 580
rect 976 570 977 580
rect 468 523 469 533
rect 471 523 472 533
rect 1332 533 1333 543
rect 1335 533 1336 543
rect 376 501 377 511
rect 380 501 382 511
rect 395 501 396 511
rect 398 501 399 511
rect 407 501 408 511
rect 410 501 411 511
rect 419 501 420 511
rect 422 501 423 511
rect 431 501 432 511
rect 434 501 435 511
rect 443 501 444 511
rect 446 501 447 511
rect 1101 505 1102 525
rect 1104 505 1114 525
rect 1116 505 1117 525
rect 1125 505 1126 525
rect 1128 505 1138 525
rect 1140 505 1141 525
rect 1367 533 1368 543
rect 1370 533 1380 543
rect 1382 533 1383 543
rect 1400 533 1401 543
rect 1403 533 1413 543
rect 1415 533 1416 543
rect 1432 533 1433 543
rect 1435 533 1436 543
rect -566 441 -565 451
rect -563 441 -553 451
rect -551 441 -550 451
rect -533 441 -532 451
rect -530 441 -520 451
rect -518 441 -517 451
rect -501 441 -500 451
rect -498 441 -497 451
rect -62 446 -61 466
rect -59 446 -49 466
rect -47 446 -46 466
rect -25 462 -24 472
rect -22 462 -21 472
rect 975 454 976 464
rect 978 454 979 464
rect -305 400 -304 420
rect -302 400 -292 420
rect -290 400 -289 420
rect -281 400 -280 420
rect -278 400 -268 420
rect -266 400 -265 420
rect -438 388 -437 398
rect -435 388 -434 398
rect 24 345 25 365
rect 27 345 37 365
rect 39 345 40 365
rect 61 361 62 371
rect 64 361 65 371
rect 129 325 130 345
rect 132 325 142 345
rect 144 325 145 345
rect 166 341 167 351
rect 169 341 170 351
rect 255 266 256 286
rect 258 266 268 286
rect 270 266 271 286
rect 292 282 293 292
rect 295 282 296 292
rect -437 200 -436 210
rect -434 200 -433 210
rect -599 143 -598 153
rect -596 143 -595 153
rect -564 143 -563 153
rect -561 143 -551 153
rect -549 143 -548 153
rect -531 143 -530 153
rect -528 143 -518 153
rect -516 143 -515 153
rect -499 143 -498 153
rect -496 143 -495 153
rect 973 170 974 180
rect 976 170 977 180
rect -382 116 -381 136
rect -379 116 -369 136
rect -367 116 -366 136
rect -345 132 -344 142
rect -342 132 -341 142
rect -102 133 -101 153
rect -99 133 -89 153
rect -87 133 -86 153
rect -65 149 -64 159
rect -62 149 -61 159
rect -601 41 -600 51
rect -598 41 -597 51
rect 1332 133 1333 143
rect 1335 133 1336 143
rect 440 111 441 121
rect 443 111 444 121
rect 367 99 368 109
rect 370 99 371 109
rect 379 99 380 109
rect 382 99 383 109
rect 391 99 392 109
rect 394 99 395 109
rect 403 99 404 109
rect 406 99 407 109
rect 415 99 416 109
rect 418 99 419 109
rect 1101 105 1102 125
rect 1104 105 1114 125
rect 1116 105 1117 125
rect 1125 105 1126 125
rect 1128 105 1138 125
rect 1140 105 1141 125
rect 1367 133 1368 143
rect 1370 133 1380 143
rect 1382 133 1383 143
rect 1400 133 1401 143
rect 1403 133 1413 143
rect 1415 133 1416 143
rect 1432 133 1433 143
rect 1435 133 1436 143
rect -566 41 -565 51
rect -563 41 -553 51
rect -551 41 -550 51
rect -533 41 -532 51
rect -530 41 -520 51
rect -518 41 -517 51
rect -501 41 -500 51
rect -498 41 -497 51
rect 17 52 18 72
rect 20 52 30 72
rect 32 52 33 72
rect 54 68 55 78
rect 57 68 58 78
rect 975 54 976 64
rect 978 54 979 64
rect -305 0 -304 20
rect -302 0 -292 20
rect -290 0 -289 20
rect -281 0 -280 20
rect -278 0 -268 20
rect -266 0 -265 20
rect -438 -12 -437 -2
rect -435 -12 -434 -2
rect 132 -44 133 -24
rect 135 -44 145 -24
rect 147 -44 148 -24
rect 169 -28 170 -18
rect 172 -28 173 -18
rect 260 -131 261 -111
rect 263 -131 273 -111
rect 275 -131 276 -111
rect 297 -115 298 -105
rect 300 -115 301 -105
rect -438 -247 -437 -237
rect -435 -247 -434 -237
rect -601 -304 -600 -294
rect -598 -304 -597 -294
rect -566 -304 -565 -294
rect -563 -304 -553 -294
rect -551 -304 -550 -294
rect -533 -304 -532 -294
rect -530 -304 -520 -294
rect -518 -304 -517 -294
rect -501 -304 -500 -294
rect -498 -304 -497 -294
rect -383 -331 -382 -311
rect -380 -331 -370 -311
rect -368 -331 -367 -311
rect -346 -315 -345 -305
rect -343 -315 -342 -305
rect -105 -312 -104 -292
rect -102 -312 -92 -292
rect -90 -312 -89 -292
rect -68 -296 -67 -286
rect -65 -296 -64 -286
rect 964 -288 965 -278
rect 967 -288 968 -278
rect 374 -312 375 -302
rect 377 -312 378 -302
rect 313 -332 314 -322
rect 316 -332 317 -322
rect 325 -332 326 -322
rect 328 -332 329 -322
rect 337 -332 338 -322
rect 340 -332 341 -322
rect 349 -332 350 -322
rect 352 -332 353 -322
rect 1329 -328 1330 -318
rect 1332 -328 1333 -318
rect -602 -406 -601 -396
rect -599 -406 -598 -396
rect 1092 -353 1093 -333
rect 1095 -353 1105 -333
rect 1107 -353 1108 -333
rect 1116 -353 1117 -333
rect 1119 -353 1129 -333
rect 1131 -353 1132 -333
rect 1364 -328 1365 -318
rect 1367 -328 1377 -318
rect 1379 -328 1380 -318
rect 1397 -328 1398 -318
rect 1400 -328 1410 -318
rect 1412 -328 1413 -318
rect 1429 -328 1430 -318
rect 1432 -328 1433 -318
rect -567 -406 -566 -396
rect -564 -406 -554 -396
rect -552 -406 -551 -396
rect -534 -406 -533 -396
rect -531 -406 -521 -396
rect -519 -406 -518 -396
rect -502 -406 -501 -396
rect -499 -406 -498 -396
rect 26 -384 27 -364
rect 29 -384 39 -364
rect 41 -384 42 -364
rect 63 -368 64 -358
rect 66 -368 67 -358
rect 966 -404 967 -394
rect 969 -404 970 -394
rect -306 -447 -305 -427
rect -303 -447 -293 -427
rect -291 -447 -290 -427
rect -282 -447 -281 -427
rect -279 -447 -269 -427
rect -267 -447 -266 -427
rect -439 -459 -438 -449
rect -436 -459 -435 -449
rect 169 -467 170 -447
rect 172 -467 182 -447
rect 184 -467 185 -447
rect 206 -451 207 -441
rect 209 -451 210 -441
rect -436 -708 -435 -698
rect -433 -708 -432 -698
rect -603 -765 -602 -755
rect -600 -765 -599 -755
rect -568 -765 -567 -755
rect -565 -765 -555 -755
rect -553 -765 -552 -755
rect -535 -765 -534 -755
rect -532 -765 -522 -755
rect -520 -765 -519 -755
rect -503 -765 -502 -755
rect -500 -765 -499 -755
rect -381 -792 -380 -772
rect -378 -792 -368 -772
rect -366 -792 -365 -772
rect -344 -776 -343 -766
rect -341 -776 -340 -766
rect 186 -779 187 -769
rect 189 -779 190 -769
rect -601 -868 -600 -858
rect -598 -868 -597 -858
rect -84 -821 -83 -801
rect -81 -821 -71 -801
rect -69 -821 -68 -801
rect -47 -805 -46 -795
rect -44 -805 -43 -795
rect 137 -799 138 -789
rect 140 -799 141 -789
rect 149 -799 150 -789
rect 152 -799 153 -789
rect 161 -799 162 -789
rect 164 -799 165 -789
rect 926 -797 927 -787
rect 929 -797 930 -787
rect -566 -868 -565 -858
rect -563 -868 -553 -858
rect -551 -868 -550 -858
rect -533 -868 -532 -858
rect -530 -868 -520 -858
rect -518 -868 -517 -858
rect -501 -868 -500 -858
rect -498 -868 -497 -858
rect 1054 -862 1055 -842
rect 1057 -862 1067 -842
rect 1069 -862 1070 -842
rect 1078 -862 1079 -842
rect 1081 -862 1091 -842
rect 1093 -862 1094 -842
rect -304 -908 -303 -888
rect -301 -908 -291 -888
rect -289 -908 -288 -888
rect -280 -908 -279 -888
rect -277 -908 -267 -888
rect -265 -908 -264 -888
rect 1332 -864 1333 -854
rect 1335 -864 1336 -854
rect 1367 -864 1368 -854
rect 1370 -864 1380 -854
rect 1382 -864 1383 -854
rect 1400 -864 1401 -854
rect 1403 -864 1413 -854
rect 1415 -864 1416 -854
rect 1432 -864 1433 -854
rect 1435 -864 1436 -854
rect -437 -920 -436 -910
rect -434 -920 -433 -910
rect 17 -913 18 -893
rect 20 -913 30 -893
rect 32 -913 33 -893
rect 54 -897 55 -887
rect 57 -897 58 -887
rect 928 -913 929 -903
rect 931 -913 932 -903
rect -683 -1072 -682 -1062
rect -680 -1072 -679 -1062
rect -648 -1072 -647 -1062
rect -645 -1072 -635 -1062
rect -633 -1072 -632 -1062
rect -615 -1072 -614 -1062
rect -612 -1072 -602 -1062
rect -600 -1072 -599 -1062
rect -583 -1072 -582 -1062
rect -580 -1072 -579 -1062
rect -435 -1162 -434 -1152
rect -432 -1162 -431 -1152
rect -601 -1215 -600 -1205
rect -598 -1215 -597 -1205
rect -566 -1215 -565 -1205
rect -563 -1215 -553 -1205
rect -551 -1215 -550 -1205
rect -533 -1215 -532 -1205
rect -530 -1215 -520 -1205
rect -518 -1215 -517 -1205
rect -501 -1215 -500 -1205
rect -498 -1215 -497 -1205
rect -380 -1246 -379 -1226
rect -377 -1246 -367 -1226
rect -365 -1246 -364 -1226
rect -343 -1230 -342 -1220
rect -340 -1230 -339 -1220
rect -111 -1228 -110 -1208
rect -108 -1228 -98 -1208
rect -96 -1228 -95 -1208
rect -74 -1212 -73 -1202
rect -71 -1212 -70 -1202
rect 902 -1220 903 -1210
rect 905 -1220 906 -1210
rect -600 -1325 -599 -1315
rect -597 -1325 -596 -1315
rect -565 -1325 -564 -1315
rect -562 -1325 -552 -1315
rect -550 -1325 -549 -1315
rect -532 -1325 -531 -1315
rect -529 -1325 -519 -1315
rect -517 -1325 -516 -1315
rect -500 -1325 -499 -1315
rect -497 -1325 -496 -1315
rect 1030 -1285 1031 -1265
rect 1033 -1285 1043 -1265
rect 1045 -1285 1046 -1265
rect 1054 -1285 1055 -1265
rect 1057 -1285 1067 -1265
rect 1069 -1285 1070 -1265
rect 1324 -1274 1325 -1264
rect 1327 -1274 1328 -1264
rect 5 -1314 6 -1304
rect 8 -1314 9 -1304
rect 17 -1314 18 -1304
rect 20 -1314 21 -1304
rect 42 -1308 43 -1298
rect 45 -1308 46 -1298
rect 1359 -1274 1360 -1264
rect 1362 -1274 1372 -1264
rect 1374 -1274 1375 -1264
rect 1392 -1274 1393 -1264
rect 1395 -1274 1405 -1264
rect 1407 -1274 1408 -1264
rect 1424 -1274 1425 -1264
rect 1427 -1274 1428 -1264
rect 904 -1336 905 -1326
rect 907 -1336 908 -1326
rect -303 -1362 -302 -1342
rect -300 -1362 -290 -1342
rect -288 -1362 -287 -1342
rect -279 -1362 -278 -1342
rect -276 -1362 -266 -1342
rect -264 -1362 -263 -1342
rect -436 -1374 -435 -1364
rect -433 -1374 -432 -1364
<< pdiffusion >>
rect 1338 950 1339 970
rect 1341 950 1351 970
rect 1353 950 1354 970
rect 1373 950 1374 970
rect 1376 950 1377 970
rect 1406 950 1407 970
rect 1409 950 1410 970
rect 1438 950 1439 970
rect 1441 950 1442 970
rect -437 630 -436 650
rect -434 630 -433 650
rect -599 574 -598 594
rect -596 574 -586 594
rect -584 574 -583 594
rect -564 574 -563 594
rect -561 574 -560 594
rect -531 574 -530 594
rect -528 574 -527 594
rect -499 574 -498 594
rect -496 574 -495 594
rect -135 585 -134 605
rect -132 585 -131 605
rect -123 585 -122 605
rect -120 585 -119 605
rect -98 586 -97 606
rect -95 586 -94 606
rect -382 561 -381 581
rect -379 561 -378 581
rect -370 561 -369 581
rect -367 561 -366 581
rect -345 562 -344 582
rect -342 562 -341 582
rect 376 573 377 699
rect 380 573 396 699
rect 398 573 408 699
rect 410 573 420 699
rect 422 573 432 699
rect 434 573 444 699
rect 446 573 447 699
rect 973 600 974 620
rect 976 600 977 620
rect -601 472 -600 492
rect -598 472 -588 492
rect -586 472 -585 492
rect -566 472 -565 492
rect -563 472 -562 492
rect -533 472 -532 492
rect -530 472 -529 492
rect -501 472 -500 492
rect -498 472 -497 492
rect -305 465 -304 505
rect -302 465 -292 505
rect -290 465 -289 505
rect -281 465 -280 505
rect -278 465 -268 505
rect -266 465 -265 505
rect -62 491 -61 511
rect -59 491 -58 511
rect -50 491 -49 511
rect -47 491 -46 511
rect -25 492 -24 512
rect -22 492 -21 512
rect 468 553 469 573
rect 471 553 472 573
rect 1101 570 1102 610
rect 1104 570 1114 610
rect 1116 570 1117 610
rect 1125 570 1126 610
rect 1128 570 1138 610
rect 1140 570 1141 610
rect 1332 564 1333 584
rect 1335 564 1345 584
rect 1347 564 1348 584
rect 1367 564 1368 584
rect 1370 564 1371 584
rect 1400 564 1401 584
rect 1403 564 1404 584
rect 1432 564 1433 584
rect 1435 564 1436 584
rect 975 484 976 504
rect 978 484 979 504
rect -438 418 -437 438
rect -435 418 -434 438
rect 24 390 25 410
rect 27 390 28 410
rect 36 390 37 410
rect 39 390 40 410
rect 61 391 62 411
rect 64 391 65 411
rect 129 370 130 390
rect 132 370 133 390
rect 141 370 142 390
rect 144 370 145 390
rect 166 371 167 391
rect 169 371 170 391
rect 255 311 256 331
rect 258 311 259 331
rect 267 311 268 331
rect 270 311 271 331
rect 292 312 293 332
rect 295 312 296 332
rect -437 230 -436 250
rect -434 230 -433 250
rect -599 174 -598 194
rect -596 174 -586 194
rect -584 174 -583 194
rect -564 174 -563 194
rect -561 174 -560 194
rect -531 174 -530 194
rect -528 174 -527 194
rect -499 174 -498 194
rect -496 174 -495 194
rect -382 161 -381 181
rect -379 161 -378 181
rect -370 161 -369 181
rect -367 161 -366 181
rect -345 162 -344 182
rect -342 162 -341 182
rect -102 178 -101 198
rect -99 178 -98 198
rect -90 178 -89 198
rect -87 178 -86 198
rect -65 179 -64 199
rect -62 179 -61 199
rect 367 161 368 261
rect 370 161 380 261
rect 382 161 392 261
rect 394 161 404 261
rect 406 161 416 261
rect 418 161 419 261
rect 973 200 974 220
rect 976 200 977 220
rect 1101 170 1102 210
rect 1104 170 1114 210
rect 1116 170 1117 210
rect 1125 170 1126 210
rect 1128 170 1138 210
rect 1140 170 1141 210
rect -601 72 -600 92
rect -598 72 -588 92
rect -586 72 -585 92
rect -566 72 -565 92
rect -563 72 -562 92
rect -533 72 -532 92
rect -530 72 -529 92
rect -501 72 -500 92
rect -498 72 -497 92
rect -305 65 -304 105
rect -302 65 -292 105
rect -290 65 -289 105
rect -281 65 -280 105
rect -278 65 -268 105
rect -266 65 -265 105
rect 17 97 18 117
rect 20 97 21 117
rect 29 97 30 117
rect 32 97 33 117
rect 54 98 55 118
rect 57 98 58 118
rect 440 141 441 161
rect 443 141 444 161
rect 1332 164 1333 184
rect 1335 164 1345 184
rect 1347 164 1348 184
rect 1367 164 1368 184
rect 1370 164 1371 184
rect 1400 164 1401 184
rect 1403 164 1404 184
rect 1432 164 1433 184
rect 1435 164 1436 184
rect 975 84 976 104
rect 978 84 979 104
rect -438 18 -437 38
rect -435 18 -434 38
rect 132 1 133 21
rect 135 1 136 21
rect 144 1 145 21
rect 147 1 148 21
rect 169 2 170 22
rect 172 2 173 22
rect 260 -86 261 -66
rect 263 -86 264 -66
rect 272 -86 273 -66
rect 275 -86 276 -66
rect 297 -85 298 -65
rect 300 -85 301 -65
rect -438 -217 -437 -197
rect -435 -217 -434 -197
rect -601 -273 -600 -253
rect -598 -273 -588 -253
rect -586 -273 -585 -253
rect -566 -273 -565 -253
rect -563 -273 -562 -253
rect -533 -273 -532 -253
rect -530 -273 -529 -253
rect -501 -273 -500 -253
rect -498 -273 -497 -253
rect -383 -286 -382 -266
rect -380 -286 -379 -266
rect -371 -286 -370 -266
rect -368 -286 -367 -266
rect -346 -285 -345 -265
rect -343 -285 -342 -265
rect -105 -267 -104 -247
rect -102 -267 -101 -247
rect -93 -267 -92 -247
rect -90 -267 -89 -247
rect -68 -266 -67 -246
rect -65 -266 -64 -246
rect 313 -283 314 -203
rect 316 -283 326 -203
rect 328 -283 338 -203
rect 340 -283 350 -203
rect 352 -283 353 -203
rect 964 -258 965 -238
rect 967 -258 968 -238
rect 374 -282 375 -262
rect 377 -282 378 -262
rect 26 -339 27 -319
rect 29 -339 30 -319
rect 38 -339 39 -319
rect 41 -339 42 -319
rect 63 -338 64 -318
rect 66 -338 67 -318
rect 1092 -288 1093 -248
rect 1095 -288 1105 -248
rect 1107 -288 1108 -248
rect 1116 -288 1117 -248
rect 1119 -288 1129 -248
rect 1131 -288 1132 -248
rect 1329 -297 1330 -277
rect 1332 -297 1342 -277
rect 1344 -297 1345 -277
rect 1364 -297 1365 -277
rect 1367 -297 1368 -277
rect 1397 -297 1398 -277
rect 1400 -297 1401 -277
rect 1429 -297 1430 -277
rect 1432 -297 1433 -277
rect -602 -375 -601 -355
rect -599 -375 -589 -355
rect -587 -375 -586 -355
rect -567 -375 -566 -355
rect -564 -375 -563 -355
rect -534 -375 -533 -355
rect -531 -375 -530 -355
rect -502 -375 -501 -355
rect -499 -375 -498 -355
rect -306 -382 -305 -342
rect -303 -382 -293 -342
rect -291 -382 -290 -342
rect -282 -382 -281 -342
rect -279 -382 -269 -342
rect -267 -382 -266 -342
rect 966 -374 967 -354
rect 969 -374 970 -354
rect -439 -429 -438 -409
rect -436 -429 -435 -409
rect 169 -422 170 -402
rect 172 -422 173 -402
rect 181 -422 182 -402
rect 184 -422 185 -402
rect 206 -421 207 -401
rect 209 -421 210 -401
rect -436 -678 -435 -658
rect -433 -678 -432 -658
rect -603 -734 -602 -714
rect -600 -734 -590 -714
rect -588 -734 -587 -714
rect -568 -734 -567 -714
rect -565 -734 -564 -714
rect -535 -734 -534 -714
rect -532 -734 -531 -714
rect -503 -734 -502 -714
rect -500 -734 -499 -714
rect -381 -747 -380 -727
rect -378 -747 -377 -727
rect -369 -747 -368 -727
rect -366 -747 -365 -727
rect -344 -746 -343 -726
rect -341 -746 -340 -726
rect 137 -753 138 -693
rect 140 -753 150 -693
rect 152 -753 162 -693
rect 164 -753 165 -693
rect 186 -749 187 -729
rect 189 -749 190 -729
rect -84 -776 -83 -756
rect -81 -776 -80 -756
rect -72 -776 -71 -756
rect -69 -776 -68 -756
rect -47 -775 -46 -755
rect -44 -775 -43 -755
rect 926 -767 927 -747
rect 929 -767 930 -747
rect -601 -837 -600 -817
rect -598 -837 -588 -817
rect -586 -837 -585 -817
rect -566 -837 -565 -817
rect -563 -837 -562 -817
rect -533 -837 -532 -817
rect -530 -837 -529 -817
rect -501 -837 -500 -817
rect -498 -837 -497 -817
rect -304 -843 -303 -803
rect -301 -843 -291 -803
rect -289 -843 -288 -803
rect -280 -843 -279 -803
rect -277 -843 -267 -803
rect -265 -843 -264 -803
rect 1054 -797 1055 -757
rect 1057 -797 1067 -757
rect 1069 -797 1070 -757
rect 1078 -797 1079 -757
rect 1081 -797 1091 -757
rect 1093 -797 1094 -757
rect 1332 -833 1333 -813
rect 1335 -833 1345 -813
rect 1347 -833 1348 -813
rect 1367 -833 1368 -813
rect 1370 -833 1371 -813
rect 1400 -833 1401 -813
rect 1403 -833 1404 -813
rect 1432 -833 1433 -813
rect 1435 -833 1436 -813
rect 17 -868 18 -848
rect 20 -868 21 -848
rect 29 -868 30 -848
rect 32 -868 33 -848
rect 54 -867 55 -847
rect 57 -867 58 -847
rect -437 -890 -436 -870
rect -434 -890 -433 -870
rect 928 -883 929 -863
rect 931 -883 932 -863
rect -683 -1041 -682 -1021
rect -680 -1041 -670 -1021
rect -668 -1041 -667 -1021
rect -648 -1041 -647 -1021
rect -645 -1041 -644 -1021
rect -615 -1041 -614 -1021
rect -612 -1041 -611 -1021
rect -583 -1041 -582 -1021
rect -580 -1041 -579 -1021
rect -435 -1132 -434 -1112
rect -432 -1132 -431 -1112
rect -601 -1184 -600 -1164
rect -598 -1184 -588 -1164
rect -586 -1184 -585 -1164
rect -566 -1184 -565 -1164
rect -563 -1184 -562 -1164
rect -533 -1184 -532 -1164
rect -530 -1184 -529 -1164
rect -501 -1184 -500 -1164
rect -498 -1184 -497 -1164
rect -380 -1201 -379 -1181
rect -377 -1201 -376 -1181
rect -368 -1201 -367 -1181
rect -365 -1201 -364 -1181
rect -343 -1200 -342 -1180
rect -340 -1200 -339 -1180
rect -111 -1183 -110 -1163
rect -108 -1183 -107 -1163
rect -99 -1183 -98 -1163
rect -96 -1183 -95 -1163
rect -74 -1182 -73 -1162
rect -71 -1182 -70 -1162
rect 902 -1190 903 -1170
rect 905 -1190 906 -1170
rect 1030 -1220 1031 -1180
rect 1033 -1220 1043 -1180
rect 1045 -1220 1046 -1180
rect 1054 -1220 1055 -1180
rect 1057 -1220 1067 -1180
rect 1069 -1220 1070 -1180
rect -600 -1294 -599 -1274
rect -597 -1294 -587 -1274
rect -585 -1294 -584 -1274
rect -565 -1294 -564 -1274
rect -562 -1294 -561 -1274
rect -532 -1294 -531 -1274
rect -529 -1294 -528 -1274
rect -500 -1294 -499 -1274
rect -497 -1294 -496 -1274
rect -303 -1297 -302 -1257
rect -300 -1297 -290 -1257
rect -288 -1297 -287 -1257
rect -279 -1297 -278 -1257
rect -276 -1297 -266 -1257
rect -264 -1297 -263 -1257
rect 5 -1280 6 -1240
rect 8 -1280 18 -1240
rect 20 -1280 21 -1240
rect 1324 -1243 1325 -1223
rect 1327 -1243 1337 -1223
rect 1339 -1243 1340 -1223
rect 1359 -1243 1360 -1223
rect 1362 -1243 1363 -1223
rect 1392 -1243 1393 -1223
rect 1395 -1243 1396 -1223
rect 1424 -1243 1425 -1223
rect 1427 -1243 1428 -1223
rect 42 -1278 43 -1258
rect 45 -1278 46 -1258
rect 904 -1306 905 -1286
rect 907 -1306 908 -1286
rect -436 -1344 -435 -1324
rect -433 -1344 -432 -1324
<< ndcontact >>
rect 1334 919 1338 929
rect 1342 919 1346 929
rect 1369 919 1373 929
rect 1389 919 1393 929
rect 1402 919 1406 929
rect 1422 919 1426 929
rect 1434 919 1438 929
rect 1442 919 1446 929
rect -441 600 -437 610
rect -433 600 -429 610
rect -603 543 -599 553
rect -595 543 -591 553
rect -568 543 -564 553
rect -548 543 -544 553
rect -535 543 -531 553
rect -515 543 -511 553
rect -503 543 -499 553
rect -495 543 -491 553
rect -386 516 -382 536
rect -366 516 -362 536
rect -349 532 -345 542
rect -341 532 -337 542
rect -139 540 -135 560
rect -119 540 -115 560
rect -102 556 -98 566
rect -94 556 -90 566
rect -139 531 -135 535
rect -129 531 -125 535
rect -119 531 -115 535
rect -97 531 -93 535
rect -386 507 -382 511
rect -376 507 -372 511
rect -366 507 -362 511
rect -344 507 -340 511
rect -605 441 -601 451
rect -597 441 -593 451
rect 969 570 973 580
rect 977 570 981 580
rect 464 523 468 533
rect 472 523 476 533
rect 1328 533 1332 543
rect 1336 533 1340 543
rect 372 501 376 511
rect 382 501 395 511
rect 399 501 407 511
rect 411 501 419 511
rect 423 501 431 511
rect 435 501 443 511
rect 447 501 451 511
rect 1097 505 1101 525
rect 1117 505 1125 525
rect 1141 505 1145 525
rect 1363 533 1367 543
rect 1383 533 1387 543
rect 1396 533 1400 543
rect 1416 533 1420 543
rect 1428 533 1432 543
rect 1436 533 1440 543
rect -570 441 -566 451
rect -550 441 -546 451
rect -537 441 -533 451
rect -517 441 -513 451
rect -505 441 -501 451
rect -497 441 -493 451
rect -66 446 -62 466
rect -46 446 -42 466
rect -29 462 -25 472
rect -21 462 -17 472
rect 971 454 975 464
rect 979 454 983 464
rect -66 437 -62 441
rect -56 437 -52 441
rect -46 437 -42 441
rect -24 437 -20 441
rect -309 400 -305 420
rect -289 400 -281 420
rect -265 400 -261 420
rect -442 388 -438 398
rect -434 388 -430 398
rect 20 345 24 365
rect 40 345 44 365
rect 57 361 61 371
rect 65 361 69 371
rect 20 336 24 340
rect 30 336 34 340
rect 40 336 44 340
rect 62 336 66 340
rect 125 325 129 345
rect 145 325 149 345
rect 162 341 166 351
rect 170 341 174 351
rect 125 316 129 320
rect 135 316 139 320
rect 145 316 149 320
rect 167 316 171 320
rect 251 266 255 286
rect 271 266 275 286
rect 288 282 292 292
rect 296 282 300 292
rect 251 257 255 261
rect 261 257 265 261
rect 271 257 275 261
rect 293 257 297 261
rect -441 200 -437 210
rect -433 200 -429 210
rect -603 143 -599 153
rect -595 143 -591 153
rect -568 143 -564 153
rect -548 143 -544 153
rect -535 143 -531 153
rect -515 143 -511 153
rect -503 143 -499 153
rect -495 143 -491 153
rect 969 170 973 180
rect 977 170 981 180
rect -386 116 -382 136
rect -366 116 -362 136
rect -349 132 -345 142
rect -341 132 -337 142
rect -106 133 -102 153
rect -86 133 -82 153
rect -69 149 -65 159
rect -61 149 -57 159
rect -106 124 -102 128
rect -96 124 -92 128
rect -86 124 -82 128
rect -64 124 -60 128
rect -386 107 -382 111
rect -376 107 -372 111
rect -366 107 -362 111
rect -344 107 -340 111
rect -605 41 -601 51
rect -597 41 -593 51
rect 1328 133 1332 143
rect 1336 133 1340 143
rect 436 111 440 121
rect 444 111 448 121
rect 363 99 367 109
rect 371 99 379 109
rect 383 99 391 109
rect 395 99 403 109
rect 407 99 415 109
rect 419 99 423 109
rect 1097 105 1101 125
rect 1117 105 1125 125
rect 1141 105 1145 125
rect 1363 133 1367 143
rect 1383 133 1387 143
rect 1396 133 1400 143
rect 1416 133 1420 143
rect 1428 133 1432 143
rect 1436 133 1440 143
rect -570 41 -566 51
rect -550 41 -546 51
rect -537 41 -533 51
rect -517 41 -513 51
rect -505 41 -501 51
rect -497 41 -493 51
rect 13 52 17 72
rect 33 52 37 72
rect 50 68 54 78
rect 58 68 62 78
rect 971 54 975 64
rect 979 54 983 64
rect 13 43 17 47
rect 23 43 27 47
rect 33 43 37 47
rect 55 43 59 47
rect -309 0 -305 20
rect -289 0 -281 20
rect -265 0 -261 20
rect -442 -12 -438 -2
rect -434 -12 -430 -2
rect 128 -44 132 -24
rect 148 -44 152 -24
rect 165 -28 169 -18
rect 173 -28 177 -18
rect 128 -53 132 -49
rect 138 -53 142 -49
rect 148 -53 152 -49
rect 170 -53 174 -49
rect 256 -131 260 -111
rect 276 -131 280 -111
rect 293 -115 297 -105
rect 301 -115 305 -105
rect 256 -140 260 -136
rect 266 -140 270 -136
rect 276 -140 280 -136
rect 298 -140 302 -136
rect -442 -247 -438 -237
rect -434 -247 -430 -237
rect -605 -304 -601 -294
rect -597 -304 -593 -294
rect -570 -304 -566 -294
rect -550 -304 -546 -294
rect -537 -304 -533 -294
rect -517 -304 -513 -294
rect -505 -304 -501 -294
rect -497 -304 -493 -294
rect -387 -331 -383 -311
rect -367 -331 -363 -311
rect -350 -315 -346 -305
rect -342 -315 -338 -305
rect -109 -312 -105 -292
rect -89 -312 -85 -292
rect -72 -296 -68 -286
rect -64 -296 -60 -286
rect -109 -321 -105 -317
rect -99 -321 -95 -317
rect -89 -321 -85 -317
rect -67 -321 -63 -317
rect -387 -340 -383 -336
rect -377 -340 -373 -336
rect -367 -340 -363 -336
rect -345 -340 -341 -336
rect 960 -288 964 -278
rect 968 -288 972 -278
rect 370 -312 374 -302
rect 378 -312 382 -302
rect 309 -332 313 -322
rect 317 -332 325 -322
rect 329 -332 337 -322
rect 341 -332 349 -322
rect 353 -332 357 -322
rect 1325 -328 1329 -318
rect 1333 -328 1337 -318
rect -606 -406 -602 -396
rect -598 -406 -594 -396
rect 1088 -353 1092 -333
rect 1108 -353 1116 -333
rect 1132 -353 1136 -333
rect 1360 -328 1364 -318
rect 1380 -328 1384 -318
rect 1393 -328 1397 -318
rect 1413 -328 1417 -318
rect 1425 -328 1429 -318
rect 1433 -328 1437 -318
rect -571 -406 -567 -396
rect -551 -406 -547 -396
rect -538 -406 -534 -396
rect -518 -406 -514 -396
rect -506 -406 -502 -396
rect -498 -406 -494 -396
rect 22 -384 26 -364
rect 42 -384 46 -364
rect 59 -368 63 -358
rect 67 -368 71 -358
rect 22 -393 26 -389
rect 32 -393 36 -389
rect 42 -393 46 -389
rect 64 -393 68 -389
rect 962 -404 966 -394
rect 970 -404 974 -394
rect -310 -447 -306 -427
rect -290 -447 -282 -427
rect -266 -447 -262 -427
rect -443 -459 -439 -449
rect -435 -459 -431 -449
rect 165 -467 169 -447
rect 185 -467 189 -447
rect 202 -451 206 -441
rect 210 -451 214 -441
rect 165 -476 169 -472
rect 175 -476 179 -472
rect 185 -476 189 -472
rect 207 -476 211 -472
rect -440 -708 -436 -698
rect -432 -708 -428 -698
rect -607 -765 -603 -755
rect -599 -765 -595 -755
rect -572 -765 -568 -755
rect -552 -765 -548 -755
rect -539 -765 -535 -755
rect -519 -765 -515 -755
rect -507 -765 -503 -755
rect -499 -765 -495 -755
rect -385 -792 -381 -772
rect -365 -792 -361 -772
rect -348 -776 -344 -766
rect -340 -776 -336 -766
rect -385 -801 -381 -797
rect -375 -801 -371 -797
rect -365 -801 -361 -797
rect -343 -801 -339 -797
rect 182 -779 186 -769
rect 190 -779 194 -769
rect -605 -868 -601 -858
rect -597 -868 -593 -858
rect -88 -821 -84 -801
rect -68 -821 -64 -801
rect -51 -805 -47 -795
rect -43 -805 -39 -795
rect 133 -799 137 -789
rect 141 -799 149 -789
rect 153 -799 161 -789
rect 165 -799 169 -789
rect 922 -797 926 -787
rect 930 -797 934 -787
rect -88 -830 -84 -826
rect -78 -830 -74 -826
rect -68 -830 -64 -826
rect -46 -830 -42 -826
rect -570 -868 -566 -858
rect -550 -868 -546 -858
rect -537 -868 -533 -858
rect -517 -868 -513 -858
rect -505 -868 -501 -858
rect -497 -868 -493 -858
rect 1050 -862 1054 -842
rect 1070 -862 1078 -842
rect 1094 -862 1098 -842
rect -308 -908 -304 -888
rect -288 -908 -280 -888
rect -264 -908 -260 -888
rect 1328 -864 1332 -854
rect 1336 -864 1340 -854
rect 1363 -864 1367 -854
rect 1383 -864 1387 -854
rect 1396 -864 1400 -854
rect 1416 -864 1420 -854
rect 1428 -864 1432 -854
rect 1436 -864 1440 -854
rect -441 -920 -437 -910
rect -433 -920 -429 -910
rect 13 -913 17 -893
rect 33 -913 37 -893
rect 50 -897 54 -887
rect 58 -897 62 -887
rect 924 -913 928 -903
rect 932 -913 936 -903
rect 13 -922 17 -918
rect 23 -922 27 -918
rect 33 -922 37 -918
rect 55 -922 59 -918
rect -687 -1072 -683 -1062
rect -679 -1072 -675 -1062
rect -652 -1072 -648 -1062
rect -632 -1072 -628 -1062
rect -619 -1072 -615 -1062
rect -599 -1072 -595 -1062
rect -587 -1072 -583 -1062
rect -579 -1072 -575 -1062
rect -439 -1162 -435 -1152
rect -431 -1162 -427 -1152
rect -605 -1215 -601 -1205
rect -597 -1215 -593 -1205
rect -570 -1215 -566 -1205
rect -550 -1215 -546 -1205
rect -537 -1215 -533 -1205
rect -517 -1215 -513 -1205
rect -505 -1215 -501 -1205
rect -497 -1215 -493 -1205
rect -384 -1246 -380 -1226
rect -364 -1246 -360 -1226
rect -347 -1230 -343 -1220
rect -339 -1230 -335 -1220
rect -115 -1228 -111 -1208
rect -95 -1228 -91 -1208
rect -78 -1212 -74 -1202
rect -70 -1212 -66 -1202
rect 898 -1220 902 -1210
rect 906 -1220 910 -1210
rect -115 -1237 -111 -1233
rect -105 -1237 -101 -1233
rect -95 -1237 -91 -1233
rect -73 -1237 -69 -1233
rect -384 -1255 -380 -1251
rect -374 -1255 -370 -1251
rect -364 -1255 -360 -1251
rect -342 -1255 -338 -1251
rect -604 -1325 -600 -1315
rect -596 -1325 -592 -1315
rect -569 -1325 -565 -1315
rect -549 -1325 -545 -1315
rect -536 -1325 -532 -1315
rect -516 -1325 -512 -1315
rect -504 -1325 -500 -1315
rect -496 -1325 -492 -1315
rect 1026 -1285 1030 -1265
rect 1046 -1285 1054 -1265
rect 1070 -1285 1074 -1265
rect 1320 -1274 1324 -1264
rect 1328 -1274 1332 -1264
rect 1 -1314 5 -1304
rect 9 -1314 17 -1304
rect 21 -1314 25 -1304
rect 38 -1308 42 -1298
rect 46 -1308 50 -1298
rect 1355 -1274 1359 -1264
rect 1375 -1274 1379 -1264
rect 1388 -1274 1392 -1264
rect 1408 -1274 1412 -1264
rect 1420 -1274 1424 -1264
rect 1428 -1274 1432 -1264
rect 900 -1336 904 -1326
rect 908 -1336 912 -1326
rect -307 -1362 -303 -1342
rect -287 -1362 -279 -1342
rect -263 -1362 -259 -1342
rect -440 -1374 -436 -1364
rect -432 -1374 -428 -1364
<< pdcontact >>
rect 1334 950 1338 970
rect 1354 950 1358 970
rect 1369 950 1373 970
rect 1377 950 1381 970
rect 1402 950 1406 970
rect 1410 950 1414 970
rect 1434 950 1438 970
rect 1442 950 1446 970
rect -441 630 -437 650
rect -433 630 -429 650
rect -137 612 -133 616
rect -129 612 -125 616
rect -121 612 -117 616
rect -102 612 -98 616
rect -603 574 -599 594
rect -583 574 -579 594
rect -568 574 -564 594
rect -560 574 -556 594
rect -535 574 -531 594
rect -527 574 -523 594
rect -503 574 -499 594
rect -495 574 -491 594
rect -384 588 -380 592
rect -376 588 -372 592
rect -368 588 -364 592
rect -349 588 -345 592
rect -139 585 -135 605
rect -131 585 -123 605
rect -119 585 -115 605
rect -102 586 -98 606
rect -94 586 -90 606
rect -386 561 -382 581
rect -378 561 -370 581
rect -366 561 -362 581
rect -349 562 -345 582
rect -341 562 -337 582
rect 372 573 376 699
rect 447 573 451 699
rect 969 600 973 620
rect 977 600 981 620
rect -64 518 -60 522
rect -56 518 -52 522
rect -48 518 -44 522
rect -29 518 -25 522
rect -605 472 -601 492
rect -585 472 -581 492
rect -570 472 -566 492
rect -562 472 -558 492
rect -537 472 -533 492
rect -529 472 -525 492
rect -505 472 -501 492
rect -497 472 -493 492
rect -309 465 -305 505
rect -289 465 -281 505
rect -265 465 -261 505
rect -66 491 -62 511
rect -58 491 -50 511
rect -46 491 -42 511
rect -29 492 -25 512
rect -21 492 -17 512
rect 464 553 468 573
rect 472 553 476 573
rect 1097 570 1101 610
rect 1117 570 1125 610
rect 1141 570 1145 610
rect 1328 564 1332 584
rect 1348 564 1352 584
rect 1363 564 1367 584
rect 1371 564 1375 584
rect 1396 564 1400 584
rect 1404 564 1408 584
rect 1428 564 1432 584
rect 1436 564 1440 584
rect 971 484 975 504
rect 979 484 983 504
rect -442 418 -438 438
rect -434 418 -430 438
rect 22 417 26 421
rect 30 417 34 421
rect 38 417 42 421
rect 57 417 61 421
rect 20 390 24 410
rect 28 390 36 410
rect 40 390 44 410
rect 57 391 61 411
rect 65 391 69 411
rect 127 397 131 401
rect 135 397 139 401
rect 143 397 147 401
rect 162 397 166 401
rect 125 370 129 390
rect 133 370 141 390
rect 145 370 149 390
rect 162 371 166 391
rect 170 371 174 391
rect 253 338 257 342
rect 261 338 265 342
rect 269 338 273 342
rect 288 338 292 342
rect 251 311 255 331
rect 259 311 267 331
rect 271 311 275 331
rect 288 312 292 332
rect 296 312 300 332
rect -441 230 -437 250
rect -433 230 -429 250
rect -104 205 -100 209
rect -96 205 -92 209
rect -88 205 -84 209
rect -69 205 -65 209
rect -603 174 -599 194
rect -583 174 -579 194
rect -568 174 -564 194
rect -560 174 -556 194
rect -535 174 -531 194
rect -527 174 -523 194
rect -503 174 -499 194
rect -495 174 -491 194
rect -384 188 -380 192
rect -376 188 -372 192
rect -368 188 -364 192
rect -349 188 -345 192
rect -386 161 -382 181
rect -378 161 -370 181
rect -366 161 -362 181
rect -349 162 -345 182
rect -341 162 -337 182
rect -106 178 -102 198
rect -98 178 -90 198
rect -86 178 -82 198
rect -69 179 -65 199
rect -61 179 -57 199
rect 363 161 367 261
rect 419 161 423 261
rect 969 200 973 220
rect 977 200 981 220
rect 1097 170 1101 210
rect 1117 170 1125 210
rect 1141 170 1145 210
rect 15 124 19 128
rect 23 124 27 128
rect 31 124 35 128
rect 50 124 54 128
rect -605 72 -601 92
rect -585 72 -581 92
rect -570 72 -566 92
rect -562 72 -558 92
rect -537 72 -533 92
rect -529 72 -525 92
rect -505 72 -501 92
rect -497 72 -493 92
rect -309 65 -305 105
rect -289 65 -281 105
rect -265 65 -261 105
rect 13 97 17 117
rect 21 97 29 117
rect 33 97 37 117
rect 50 98 54 118
rect 58 98 62 118
rect 436 141 440 161
rect 444 141 448 161
rect 1328 164 1332 184
rect 1348 164 1352 184
rect 1363 164 1367 184
rect 1371 164 1375 184
rect 1396 164 1400 184
rect 1404 164 1408 184
rect 1428 164 1432 184
rect 1436 164 1440 184
rect 971 84 975 104
rect 979 84 983 104
rect -442 18 -438 38
rect -434 18 -430 38
rect 130 28 134 32
rect 138 28 142 32
rect 146 28 150 32
rect 165 28 169 32
rect 128 1 132 21
rect 136 1 144 21
rect 148 1 152 21
rect 165 2 169 22
rect 173 2 177 22
rect 258 -59 262 -55
rect 266 -59 270 -55
rect 274 -59 278 -55
rect 293 -59 297 -55
rect 256 -86 260 -66
rect 264 -86 272 -66
rect 276 -86 280 -66
rect 293 -85 297 -65
rect 301 -85 305 -65
rect -442 -217 -438 -197
rect -434 -217 -430 -197
rect -107 -240 -103 -236
rect -99 -240 -95 -236
rect -91 -240 -87 -236
rect -72 -240 -68 -236
rect -605 -273 -601 -253
rect -585 -273 -581 -253
rect -570 -273 -566 -253
rect -562 -273 -558 -253
rect -537 -273 -533 -253
rect -529 -273 -525 -253
rect -505 -273 -501 -253
rect -497 -273 -493 -253
rect -385 -259 -381 -255
rect -377 -259 -373 -255
rect -369 -259 -365 -255
rect -350 -259 -346 -255
rect -387 -286 -383 -266
rect -379 -286 -371 -266
rect -367 -286 -363 -266
rect -350 -285 -346 -265
rect -342 -285 -338 -265
rect -109 -267 -105 -247
rect -101 -267 -93 -247
rect -89 -267 -85 -247
rect -72 -266 -68 -246
rect -64 -266 -60 -246
rect 309 -283 313 -203
rect 353 -283 357 -203
rect 960 -258 964 -238
rect 968 -258 972 -238
rect 370 -282 374 -262
rect 378 -282 382 -262
rect 24 -312 28 -308
rect 32 -312 36 -308
rect 40 -312 44 -308
rect 59 -312 63 -308
rect 22 -339 26 -319
rect 30 -339 38 -319
rect 42 -339 46 -319
rect 59 -338 63 -318
rect 67 -338 71 -318
rect 1088 -288 1092 -248
rect 1108 -288 1116 -248
rect 1132 -288 1136 -248
rect 1325 -297 1329 -277
rect 1345 -297 1349 -277
rect 1360 -297 1364 -277
rect 1368 -297 1372 -277
rect 1393 -297 1397 -277
rect 1401 -297 1405 -277
rect 1425 -297 1429 -277
rect 1433 -297 1437 -277
rect -606 -375 -602 -355
rect -586 -375 -582 -355
rect -571 -375 -567 -355
rect -563 -375 -559 -355
rect -538 -375 -534 -355
rect -530 -375 -526 -355
rect -506 -375 -502 -355
rect -498 -375 -494 -355
rect -310 -382 -306 -342
rect -290 -382 -282 -342
rect -266 -382 -262 -342
rect 962 -374 966 -354
rect 970 -374 974 -354
rect 167 -395 171 -391
rect 175 -395 179 -391
rect 183 -395 187 -391
rect 202 -395 206 -391
rect -443 -429 -439 -409
rect -435 -429 -431 -409
rect 165 -422 169 -402
rect 173 -422 181 -402
rect 185 -422 189 -402
rect 202 -421 206 -401
rect 210 -421 214 -401
rect -440 -678 -436 -658
rect -432 -678 -428 -658
rect -607 -734 -603 -714
rect -587 -734 -583 -714
rect -572 -734 -568 -714
rect -564 -734 -560 -714
rect -539 -734 -535 -714
rect -531 -734 -527 -714
rect -507 -734 -503 -714
rect -499 -734 -495 -714
rect -383 -720 -379 -716
rect -375 -720 -371 -716
rect -367 -720 -363 -716
rect -348 -720 -344 -716
rect -385 -747 -381 -727
rect -377 -747 -369 -727
rect -365 -747 -361 -727
rect -348 -746 -344 -726
rect -340 -746 -336 -726
rect -86 -749 -82 -745
rect -78 -749 -74 -745
rect -70 -749 -66 -745
rect -51 -749 -47 -745
rect 133 -753 137 -693
rect 165 -753 169 -693
rect 182 -749 186 -729
rect 190 -749 194 -729
rect -88 -776 -84 -756
rect -80 -776 -72 -756
rect -68 -776 -64 -756
rect -51 -775 -47 -755
rect -43 -775 -39 -755
rect 922 -767 926 -747
rect 930 -767 934 -747
rect -605 -837 -601 -817
rect -585 -837 -581 -817
rect -570 -837 -566 -817
rect -562 -837 -558 -817
rect -537 -837 -533 -817
rect -529 -837 -525 -817
rect -505 -837 -501 -817
rect -497 -837 -493 -817
rect -308 -843 -304 -803
rect -288 -843 -280 -803
rect -264 -843 -260 -803
rect 1050 -797 1054 -757
rect 1070 -797 1078 -757
rect 1094 -797 1098 -757
rect 15 -841 19 -837
rect 23 -841 27 -837
rect 31 -841 35 -837
rect 50 -841 54 -837
rect 1328 -833 1332 -813
rect 1348 -833 1352 -813
rect 1363 -833 1367 -813
rect 1371 -833 1375 -813
rect 1396 -833 1400 -813
rect 1404 -833 1408 -813
rect 1428 -833 1432 -813
rect 1436 -833 1440 -813
rect 13 -868 17 -848
rect 21 -868 29 -848
rect 33 -868 37 -848
rect 50 -867 54 -847
rect 58 -867 62 -847
rect -441 -890 -437 -870
rect -433 -890 -429 -870
rect 924 -883 928 -863
rect 932 -883 936 -863
rect -687 -1041 -683 -1021
rect -667 -1041 -663 -1021
rect -652 -1041 -648 -1021
rect -644 -1041 -640 -1021
rect -619 -1041 -615 -1021
rect -611 -1041 -607 -1021
rect -587 -1041 -583 -1021
rect -579 -1041 -575 -1021
rect -439 -1132 -435 -1112
rect -431 -1132 -427 -1112
rect -113 -1156 -109 -1152
rect -105 -1156 -101 -1152
rect -97 -1156 -93 -1152
rect -78 -1156 -74 -1152
rect -605 -1184 -601 -1164
rect -585 -1184 -581 -1164
rect -570 -1184 -566 -1164
rect -562 -1184 -558 -1164
rect -537 -1184 -533 -1164
rect -529 -1184 -525 -1164
rect -505 -1184 -501 -1164
rect -497 -1184 -493 -1164
rect -382 -1174 -378 -1170
rect -374 -1174 -370 -1170
rect -366 -1174 -362 -1170
rect -347 -1174 -343 -1170
rect -384 -1201 -380 -1181
rect -376 -1201 -368 -1181
rect -364 -1201 -360 -1181
rect -347 -1200 -343 -1180
rect -339 -1200 -335 -1180
rect -115 -1183 -111 -1163
rect -107 -1183 -99 -1163
rect -95 -1183 -91 -1163
rect -78 -1182 -74 -1162
rect -70 -1182 -66 -1162
rect 898 -1190 902 -1170
rect 906 -1190 910 -1170
rect 1026 -1220 1030 -1180
rect 1046 -1220 1054 -1180
rect 1070 -1220 1074 -1180
rect -604 -1294 -600 -1274
rect -584 -1294 -580 -1274
rect -569 -1294 -565 -1274
rect -561 -1294 -557 -1274
rect -536 -1294 -532 -1274
rect -528 -1294 -524 -1274
rect -504 -1294 -500 -1274
rect -496 -1294 -492 -1274
rect -307 -1297 -303 -1257
rect -287 -1297 -279 -1257
rect -263 -1297 -259 -1257
rect 1 -1280 5 -1240
rect 21 -1280 25 -1240
rect 1320 -1243 1324 -1223
rect 1340 -1243 1344 -1223
rect 1355 -1243 1359 -1223
rect 1363 -1243 1367 -1223
rect 1388 -1243 1392 -1223
rect 1396 -1243 1400 -1223
rect 1420 -1243 1424 -1223
rect 1428 -1243 1432 -1223
rect 38 -1278 42 -1258
rect 46 -1278 50 -1258
rect 900 -1306 904 -1286
rect 908 -1306 912 -1286
rect -440 -1344 -436 -1324
rect -432 -1344 -428 -1324
<< psubstratepdiff >>
rect 391 492 395 496
<< nsubstratendiff >>
rect 392 705 395 709
<< psubstratepcontact >>
rect 1334 911 1338 915
rect 1369 911 1373 915
rect 1378 911 1382 915
rect 1389 911 1393 915
rect 1402 911 1406 915
rect 1412 911 1416 915
rect 1422 911 1426 915
rect 1434 911 1438 915
rect -603 535 -599 539
rect -568 535 -564 539
rect -559 535 -555 539
rect -548 535 -544 539
rect -535 535 -531 539
rect -525 535 -521 539
rect -515 535 -511 539
rect -503 535 -499 539
rect -605 433 -601 437
rect 1328 525 1332 529
rect 464 511 468 515
rect 1363 525 1367 529
rect 1372 525 1376 529
rect 1383 525 1387 529
rect 1396 525 1400 529
rect 1406 525 1410 529
rect 1416 525 1420 529
rect 1428 525 1432 529
rect 385 493 391 497
rect 401 492 405 496
rect 413 492 417 496
rect 425 492 429 496
rect 437 492 441 496
rect 447 492 451 496
rect 1097 496 1101 500
rect 1107 496 1111 500
rect 1119 496 1123 500
rect 1131 496 1135 500
rect 1141 496 1145 500
rect -570 433 -566 437
rect -561 433 -557 437
rect -550 433 -546 437
rect -537 433 -533 437
rect -527 433 -523 437
rect -517 433 -513 437
rect -505 433 -501 437
rect -309 391 -305 395
rect -299 391 -295 395
rect -287 391 -283 395
rect -275 391 -271 395
rect -265 391 -261 395
rect -603 135 -599 139
rect -568 135 -564 139
rect -559 135 -555 139
rect -548 135 -544 139
rect -535 135 -531 139
rect -525 135 -521 139
rect -515 135 -511 139
rect -503 135 -499 139
rect -605 33 -601 37
rect 1328 125 1332 129
rect 1363 125 1367 129
rect 1372 125 1376 129
rect 1383 125 1387 129
rect 1396 125 1400 129
rect 1406 125 1410 129
rect 1416 125 1420 129
rect 1428 125 1432 129
rect 436 99 440 103
rect 363 90 367 94
rect 373 90 377 94
rect 385 90 389 94
rect 397 90 401 94
rect 409 90 413 94
rect 419 90 423 94
rect 1097 96 1101 100
rect 1107 96 1111 100
rect 1119 96 1123 100
rect 1131 96 1135 100
rect 1141 96 1145 100
rect -570 33 -566 37
rect -561 33 -557 37
rect -550 33 -546 37
rect -537 33 -533 37
rect -527 33 -523 37
rect -517 33 -513 37
rect -505 33 -501 37
rect -309 -9 -305 -5
rect -299 -9 -295 -5
rect -287 -9 -283 -5
rect -275 -9 -271 -5
rect -265 -9 -261 -5
rect -605 -312 -601 -308
rect -570 -312 -566 -308
rect -561 -312 -557 -308
rect -550 -312 -546 -308
rect -537 -312 -533 -308
rect -527 -312 -523 -308
rect -517 -312 -513 -308
rect -505 -312 -501 -308
rect 370 -326 374 -322
rect -606 -414 -602 -410
rect 309 -340 313 -336
rect 319 -340 323 -336
rect 331 -340 335 -336
rect 343 -340 347 -336
rect 353 -340 357 -336
rect 1325 -336 1329 -332
rect 1360 -336 1364 -332
rect 1369 -336 1373 -332
rect 1380 -336 1384 -332
rect 1393 -336 1397 -332
rect 1403 -336 1407 -332
rect 1413 -336 1417 -332
rect 1425 -336 1429 -332
rect 1088 -362 1092 -358
rect 1098 -362 1102 -358
rect 1110 -362 1114 -358
rect 1122 -362 1126 -358
rect 1132 -362 1136 -358
rect -571 -414 -567 -410
rect -562 -414 -558 -410
rect -551 -414 -547 -410
rect -538 -414 -534 -410
rect -528 -414 -524 -410
rect -518 -414 -514 -410
rect -506 -414 -502 -410
rect -310 -456 -306 -452
rect -300 -456 -296 -452
rect -288 -456 -284 -452
rect -276 -456 -272 -452
rect -266 -456 -262 -452
rect -607 -773 -603 -769
rect -572 -773 -568 -769
rect -563 -773 -559 -769
rect -552 -773 -548 -769
rect -539 -773 -535 -769
rect -529 -773 -525 -769
rect -519 -773 -515 -769
rect -507 -773 -503 -769
rect -605 -876 -601 -872
rect 133 -809 137 -805
rect 143 -809 147 -805
rect 155 -809 159 -805
rect 165 -809 169 -805
rect -570 -876 -566 -872
rect -561 -876 -557 -872
rect -550 -876 -546 -872
rect -537 -876 -533 -872
rect -527 -876 -523 -872
rect -517 -876 -513 -872
rect -505 -876 -501 -872
rect 1050 -871 1054 -867
rect 1060 -871 1064 -867
rect 1072 -871 1076 -867
rect 1084 -871 1088 -867
rect 1094 -871 1098 -867
rect 1328 -872 1332 -868
rect 1363 -872 1367 -868
rect 1372 -872 1376 -868
rect 1383 -872 1387 -868
rect 1396 -872 1400 -868
rect 1406 -872 1410 -868
rect 1416 -872 1420 -868
rect 1428 -872 1432 -868
rect -308 -917 -304 -913
rect -298 -917 -294 -913
rect -286 -917 -282 -913
rect -274 -917 -270 -913
rect -264 -917 -260 -913
rect -687 -1080 -683 -1076
rect -652 -1080 -648 -1076
rect -643 -1080 -639 -1076
rect -632 -1080 -628 -1076
rect -619 -1080 -615 -1076
rect -609 -1080 -605 -1076
rect -599 -1080 -595 -1076
rect -587 -1080 -583 -1076
rect -605 -1223 -601 -1219
rect -570 -1223 -566 -1219
rect -561 -1223 -557 -1219
rect -550 -1223 -546 -1219
rect -537 -1223 -533 -1219
rect -527 -1223 -523 -1219
rect -517 -1223 -513 -1219
rect -505 -1223 -501 -1219
rect -604 -1333 -600 -1329
rect 1320 -1282 1324 -1278
rect 1355 -1282 1359 -1278
rect 1364 -1282 1368 -1278
rect 1375 -1282 1379 -1278
rect 1388 -1282 1392 -1278
rect 1398 -1282 1402 -1278
rect 1408 -1282 1412 -1278
rect 1420 -1282 1424 -1278
rect 1026 -1294 1030 -1290
rect 1036 -1294 1040 -1290
rect 1048 -1294 1052 -1290
rect 1060 -1294 1064 -1290
rect 1070 -1294 1074 -1290
rect 43 -1318 47 -1314
rect 1 -1324 5 -1320
rect 11 -1324 15 -1320
rect 21 -1324 25 -1320
rect -569 -1333 -565 -1329
rect -560 -1333 -556 -1329
rect -549 -1333 -545 -1329
rect -536 -1333 -532 -1329
rect -526 -1333 -522 -1329
rect -516 -1333 -512 -1329
rect -504 -1333 -500 -1329
rect -307 -1371 -303 -1367
rect -297 -1371 -293 -1367
rect -285 -1371 -281 -1367
rect -273 -1371 -269 -1367
rect -263 -1371 -259 -1367
<< nsubstratencontact >>
rect 1334 974 1338 978
rect 1344 974 1348 978
rect 1354 974 1358 978
rect 1374 974 1378 978
rect 1402 974 1406 978
rect 1434 974 1438 978
rect 384 705 392 709
rect 400 705 404 709
rect 412 705 416 709
rect 424 705 428 709
rect 436 705 440 709
rect 446 705 450 709
rect -603 598 -599 602
rect -593 598 -589 602
rect -583 598 -579 602
rect -563 598 -559 602
rect -535 598 -531 602
rect -503 598 -499 602
rect 1097 615 1101 619
rect 1107 615 1111 619
rect 1119 615 1123 619
rect 1130 615 1134 619
rect 1141 615 1145 619
rect 464 581 468 586
rect -309 510 -305 514
rect -299 510 -295 514
rect -287 510 -283 514
rect -276 510 -272 514
rect -265 510 -261 514
rect -605 496 -601 500
rect -595 496 -591 500
rect -585 496 -581 500
rect -565 496 -561 500
rect -537 496 -533 500
rect -505 496 -501 500
rect 1328 588 1332 592
rect 1338 588 1342 592
rect 1348 588 1352 592
rect 1368 588 1372 592
rect 1396 588 1400 592
rect 1428 588 1432 592
rect 363 266 367 270
rect 372 266 376 270
rect 384 266 388 270
rect 396 266 400 270
rect 408 266 412 270
rect 418 266 422 270
rect -603 198 -599 202
rect -593 198 -589 202
rect -583 198 -579 202
rect -563 198 -559 202
rect -535 198 -531 202
rect -503 198 -499 202
rect 1097 215 1101 219
rect 1107 215 1111 219
rect 1119 215 1123 219
rect 1130 215 1134 219
rect 1141 215 1145 219
rect 436 169 440 174
rect 1328 188 1332 192
rect 1338 188 1342 192
rect 1348 188 1352 192
rect 1368 188 1372 192
rect 1396 188 1400 192
rect 1428 188 1432 192
rect -309 110 -305 114
rect -299 110 -295 114
rect -287 110 -283 114
rect -276 110 -272 114
rect -265 110 -261 114
rect -605 96 -601 100
rect -595 96 -591 100
rect -585 96 -581 100
rect -565 96 -561 100
rect -537 96 -533 100
rect -505 96 -501 100
rect 309 -199 313 -195
rect 318 -199 322 -195
rect 330 -199 334 -195
rect 343 -199 347 -195
rect 353 -199 357 -195
rect -605 -249 -601 -245
rect -595 -249 -591 -245
rect -585 -249 -581 -245
rect -565 -249 -561 -245
rect -537 -249 -533 -245
rect -505 -249 -501 -245
rect 370 -256 374 -252
rect 1088 -243 1092 -239
rect 1098 -243 1102 -239
rect 1110 -243 1114 -239
rect 1121 -243 1125 -239
rect 1132 -243 1136 -239
rect -310 -337 -306 -333
rect -300 -337 -296 -333
rect -288 -337 -284 -333
rect -277 -337 -273 -333
rect -266 -337 -262 -333
rect 1325 -273 1329 -269
rect 1335 -273 1339 -269
rect 1345 -273 1349 -269
rect 1365 -273 1369 -269
rect 1393 -273 1397 -269
rect 1425 -273 1429 -269
rect -606 -351 -602 -347
rect -596 -351 -592 -347
rect -586 -351 -582 -347
rect -566 -351 -562 -347
rect -538 -351 -534 -347
rect -506 -351 -502 -347
rect 133 -689 137 -685
rect 142 -689 146 -685
rect 154 -689 158 -685
rect 165 -689 169 -685
rect -607 -710 -603 -706
rect -597 -710 -593 -706
rect -587 -710 -583 -706
rect -567 -710 -563 -706
rect -539 -710 -535 -706
rect -507 -710 -503 -706
rect -308 -798 -304 -794
rect -298 -798 -294 -794
rect -286 -798 -282 -794
rect -275 -798 -271 -794
rect -264 -798 -260 -794
rect 1050 -752 1054 -748
rect 1060 -752 1064 -748
rect 1072 -752 1076 -748
rect 1083 -752 1087 -748
rect 1094 -752 1098 -748
rect -605 -813 -601 -809
rect -595 -813 -591 -809
rect -585 -813 -581 -809
rect -565 -813 -561 -809
rect -537 -813 -533 -809
rect -505 -813 -501 -809
rect 1328 -809 1332 -805
rect 1338 -809 1342 -805
rect 1348 -809 1352 -805
rect 1368 -809 1372 -805
rect 1396 -809 1400 -805
rect 1428 -809 1432 -805
rect -687 -1017 -683 -1013
rect -677 -1017 -673 -1013
rect -667 -1017 -663 -1013
rect -647 -1017 -643 -1013
rect -619 -1017 -615 -1013
rect -587 -1017 -583 -1013
rect -605 -1160 -601 -1156
rect -595 -1160 -591 -1156
rect -585 -1160 -581 -1156
rect -565 -1160 -561 -1156
rect -537 -1160 -533 -1156
rect -505 -1160 -501 -1156
rect 1026 -1175 1030 -1171
rect 1036 -1175 1040 -1171
rect 1048 -1175 1052 -1171
rect 1059 -1175 1063 -1171
rect 1070 -1175 1074 -1171
rect 1320 -1219 1324 -1215
rect 1330 -1219 1334 -1215
rect 1340 -1219 1344 -1215
rect 1360 -1219 1364 -1215
rect 1388 -1219 1392 -1215
rect 1420 -1219 1424 -1215
rect 1 -1236 5 -1232
rect 11 -1236 15 -1232
rect 21 -1236 25 -1232
rect -307 -1252 -303 -1248
rect -297 -1252 -293 -1248
rect -285 -1252 -281 -1248
rect -274 -1252 -270 -1248
rect -263 -1252 -259 -1248
rect -604 -1270 -600 -1266
rect -594 -1270 -590 -1266
rect -584 -1270 -580 -1266
rect -564 -1270 -560 -1266
rect -536 -1270 -532 -1266
rect -504 -1270 -500 -1266
rect 38 -1251 42 -1247
<< polysilicon >>
rect 1339 970 1341 973
rect 1351 970 1353 973
rect 1374 970 1376 973
rect 1407 970 1409 973
rect 1439 970 1441 973
rect 1339 929 1341 950
rect 1339 916 1341 919
rect 1351 906 1353 950
rect 1374 929 1376 950
rect 1386 929 1388 943
rect 1407 929 1409 950
rect 1419 929 1421 932
rect 1439 929 1441 950
rect 1374 906 1376 919
rect 1386 916 1388 919
rect 1407 916 1409 919
rect 1419 906 1421 919
rect 1439 916 1441 919
rect 1351 904 1421 906
rect 377 699 380 702
rect 396 699 398 702
rect 408 699 410 702
rect 420 699 422 703
rect 432 699 434 703
rect 444 699 446 703
rect -436 650 -434 653
rect -436 610 -434 630
rect -134 605 -132 609
rect -122 605 -120 609
rect -97 606 -95 609
rect -598 594 -596 597
rect -586 594 -584 597
rect -563 594 -561 597
rect -530 594 -528 597
rect -498 594 -496 597
rect -436 595 -434 600
rect -381 581 -379 585
rect -369 581 -367 585
rect -344 582 -342 585
rect -598 553 -596 574
rect -598 540 -596 543
rect -586 530 -584 574
rect -563 553 -561 574
rect -551 553 -549 567
rect -530 553 -528 574
rect -518 553 -516 556
rect -498 553 -496 574
rect -563 530 -561 543
rect -551 540 -549 543
rect -530 540 -528 543
rect -518 530 -516 543
rect -498 540 -496 543
rect -381 536 -379 561
rect -369 536 -367 561
rect -344 542 -342 562
rect -134 560 -132 585
rect -122 560 -120 585
rect -97 566 -95 586
rect 974 620 976 623
rect 1102 610 1104 613
rect 1114 610 1116 613
rect 1126 610 1128 613
rect 1138 610 1140 613
rect 974 580 976 600
rect 469 573 471 576
rect -586 528 -516 530
rect -97 551 -95 556
rect -134 536 -132 540
rect -122 536 -120 540
rect -344 527 -342 532
rect -381 512 -379 516
rect -369 512 -367 516
rect -61 511 -59 515
rect -49 511 -47 515
rect -24 512 -22 515
rect -304 505 -302 508
rect -292 505 -290 508
rect -280 505 -278 508
rect -268 505 -266 508
rect -600 492 -598 495
rect -588 492 -586 495
rect -565 492 -563 495
rect -532 492 -530 495
rect -500 492 -498 495
rect -600 451 -598 472
rect -600 438 -598 441
rect -588 428 -586 472
rect -565 451 -563 472
rect -553 451 -551 465
rect -532 451 -530 472
rect -520 451 -518 454
rect -500 451 -498 472
rect 377 511 380 573
rect 396 511 398 573
rect 408 511 410 573
rect 420 511 422 573
rect 432 511 434 573
rect 444 511 446 573
rect 1333 584 1335 587
rect 1345 584 1347 587
rect 1368 584 1370 587
rect 1401 584 1403 587
rect 1433 584 1435 587
rect 974 565 976 570
rect 1102 558 1104 570
rect 469 533 471 553
rect 1114 551 1116 570
rect 1126 558 1128 570
rect 1138 551 1140 570
rect 1333 543 1335 564
rect 1102 525 1104 533
rect 1114 525 1116 540
rect 1126 525 1128 532
rect 1138 525 1140 541
rect 1333 530 1335 533
rect 469 518 471 523
rect 976 504 978 507
rect 1345 520 1347 564
rect 1368 543 1370 564
rect 1380 543 1382 557
rect 1401 543 1403 564
rect 1413 543 1415 546
rect 1433 543 1435 564
rect 1368 520 1370 533
rect 1380 530 1382 533
rect 1401 530 1403 533
rect 1413 520 1415 533
rect 1433 530 1435 533
rect 1345 518 1415 520
rect 377 498 380 501
rect 396 498 398 501
rect 408 498 410 501
rect 420 498 422 501
rect 432 498 434 501
rect 444 498 446 501
rect -61 466 -59 491
rect -49 466 -47 491
rect -24 472 -22 492
rect 1102 502 1104 505
rect 1114 502 1116 505
rect 1126 502 1128 505
rect 1138 502 1140 505
rect -304 453 -302 465
rect -292 446 -290 465
rect -280 453 -278 465
rect -268 446 -266 465
rect 976 464 978 484
rect -24 457 -22 462
rect 976 449 978 454
rect -61 442 -59 446
rect -49 442 -47 446
rect -565 428 -563 441
rect -553 438 -551 441
rect -532 438 -530 441
rect -520 428 -518 441
rect -500 438 -498 441
rect -437 438 -435 441
rect -588 426 -518 428
rect -304 420 -302 428
rect -292 420 -290 435
rect -280 420 -278 427
rect -268 420 -266 436
rect -437 398 -435 418
rect 25 410 27 414
rect 37 410 39 414
rect 62 411 64 414
rect -304 397 -302 400
rect -292 397 -290 400
rect -280 397 -278 400
rect -268 397 -266 400
rect -437 383 -435 388
rect 25 365 27 390
rect 37 365 39 390
rect 62 371 64 391
rect 130 390 132 394
rect 142 390 144 394
rect 167 391 169 394
rect 62 356 64 361
rect 130 345 132 370
rect 142 345 144 370
rect 167 351 169 371
rect 25 341 27 345
rect 37 341 39 345
rect 167 336 169 341
rect 256 331 258 335
rect 268 331 270 335
rect 293 332 295 335
rect 130 321 132 325
rect 142 321 144 325
rect 256 286 258 311
rect 268 286 270 311
rect 293 292 295 312
rect 293 277 295 282
rect 256 262 258 266
rect 268 262 270 266
rect 368 261 370 264
rect 380 261 382 264
rect 392 261 394 264
rect 404 261 406 264
rect 416 261 418 264
rect -436 250 -434 253
rect -436 210 -434 230
rect -598 194 -596 197
rect -586 194 -584 197
rect -563 194 -561 197
rect -530 194 -528 197
rect -498 194 -496 197
rect -436 195 -434 200
rect -101 198 -99 202
rect -89 198 -87 202
rect -64 199 -62 202
rect -381 181 -379 185
rect -369 181 -367 185
rect -344 182 -342 185
rect -598 153 -596 174
rect -598 140 -596 143
rect -586 130 -584 174
rect -563 153 -561 174
rect -551 153 -549 167
rect -530 153 -528 174
rect -518 153 -516 156
rect -498 153 -496 174
rect -563 130 -561 143
rect -551 140 -549 143
rect -530 140 -528 143
rect -518 130 -516 143
rect -498 140 -496 143
rect -381 136 -379 161
rect -369 136 -367 161
rect -344 142 -342 162
rect -101 153 -99 178
rect -89 153 -87 178
rect -64 159 -62 179
rect 974 220 976 223
rect 1102 210 1104 213
rect 1114 210 1116 213
rect 1126 210 1128 213
rect 1138 210 1140 213
rect 974 180 976 200
rect 1333 184 1335 187
rect 1345 184 1347 187
rect 1368 184 1370 187
rect 1401 184 1403 187
rect 1433 184 1435 187
rect 974 165 976 170
rect 441 161 443 164
rect -586 128 -516 130
rect -64 144 -62 149
rect -344 127 -342 132
rect -101 129 -99 133
rect -89 129 -87 133
rect 18 117 20 121
rect 30 117 32 121
rect 55 118 57 121
rect -381 112 -379 116
rect -369 112 -367 116
rect -304 105 -302 108
rect -292 105 -290 108
rect -280 105 -278 108
rect -268 105 -266 108
rect -600 92 -598 95
rect -588 92 -586 95
rect -565 92 -563 95
rect -532 92 -530 95
rect -500 92 -498 95
rect -600 51 -598 72
rect -600 38 -598 41
rect -588 28 -586 72
rect -565 51 -563 72
rect -553 51 -551 65
rect -532 51 -530 72
rect -520 51 -518 54
rect -500 51 -498 72
rect 368 109 370 161
rect 380 109 382 161
rect 392 109 394 161
rect 404 109 406 161
rect 416 109 418 161
rect 1102 158 1104 170
rect 1114 151 1116 170
rect 1126 158 1128 170
rect 1138 151 1140 170
rect 1333 143 1335 164
rect 441 121 443 141
rect 1102 125 1104 133
rect 1114 125 1116 140
rect 1126 125 1128 132
rect 1138 125 1140 141
rect 1333 130 1335 133
rect 441 106 443 111
rect 976 104 978 107
rect 1345 120 1347 164
rect 1368 143 1370 164
rect 1380 143 1382 157
rect 1401 143 1403 164
rect 1413 143 1415 146
rect 1433 143 1435 164
rect 1368 120 1370 133
rect 1380 130 1382 133
rect 1401 130 1403 133
rect 1413 120 1415 133
rect 1433 130 1435 133
rect 1345 118 1415 120
rect 18 72 20 97
rect 30 72 32 97
rect 55 78 57 98
rect 368 96 370 99
rect 380 96 382 99
rect 392 96 394 99
rect 404 96 406 99
rect 416 96 418 99
rect 1102 102 1104 105
rect 1114 102 1116 105
rect 1126 102 1128 105
rect 1138 102 1140 105
rect -304 53 -302 65
rect -292 46 -290 65
rect -280 53 -278 65
rect -268 46 -266 65
rect 55 63 57 68
rect 976 64 978 84
rect 18 48 20 52
rect 30 48 32 52
rect 976 49 978 54
rect -565 28 -563 41
rect -553 38 -551 41
rect -532 38 -530 41
rect -520 28 -518 41
rect -500 38 -498 41
rect -437 38 -435 41
rect -588 26 -518 28
rect -304 20 -302 28
rect -292 20 -290 35
rect -280 20 -278 27
rect -268 20 -266 36
rect 133 21 135 25
rect 145 21 147 25
rect 170 22 172 25
rect -437 -2 -435 18
rect -304 -3 -302 0
rect -292 -3 -290 0
rect -280 -3 -278 0
rect -268 -3 -266 0
rect -437 -17 -435 -12
rect 133 -24 135 1
rect 145 -24 147 1
rect 170 -18 172 2
rect 170 -33 172 -28
rect 133 -48 135 -44
rect 145 -48 147 -44
rect 261 -66 263 -62
rect 273 -66 275 -62
rect 298 -65 300 -62
rect 261 -111 263 -86
rect 273 -111 275 -86
rect 298 -105 300 -85
rect 298 -120 300 -115
rect 261 -135 263 -131
rect 273 -135 275 -131
rect -437 -197 -435 -194
rect 314 -203 316 -200
rect 326 -203 328 -200
rect 338 -203 340 -200
rect 350 -203 352 -200
rect -437 -237 -435 -217
rect -104 -247 -102 -243
rect -92 -247 -90 -243
rect -67 -246 -65 -243
rect -600 -253 -598 -250
rect -588 -253 -586 -250
rect -565 -253 -563 -250
rect -532 -253 -530 -250
rect -500 -253 -498 -250
rect -437 -252 -435 -247
rect -382 -266 -380 -262
rect -370 -266 -368 -262
rect -345 -265 -343 -262
rect -600 -294 -598 -273
rect -600 -307 -598 -304
rect -588 -317 -586 -273
rect -565 -294 -563 -273
rect -553 -294 -551 -280
rect -532 -294 -530 -273
rect -520 -294 -518 -291
rect -500 -294 -498 -273
rect -565 -317 -563 -304
rect -553 -307 -551 -304
rect -532 -307 -530 -304
rect -520 -317 -518 -304
rect -500 -307 -498 -304
rect -382 -311 -380 -286
rect -370 -311 -368 -286
rect -345 -305 -343 -285
rect -104 -292 -102 -267
rect -92 -292 -90 -267
rect -67 -286 -65 -266
rect 965 -238 967 -235
rect 1093 -248 1095 -245
rect 1105 -248 1107 -245
rect 1117 -248 1119 -245
rect 1129 -248 1131 -245
rect 375 -262 377 -259
rect 965 -278 967 -258
rect -588 -319 -518 -317
rect -67 -301 -65 -296
rect -345 -320 -343 -315
rect -104 -316 -102 -312
rect -92 -316 -90 -312
rect 27 -319 29 -315
rect 39 -319 41 -315
rect 64 -318 66 -315
rect -382 -335 -380 -331
rect -370 -335 -368 -331
rect 314 -322 316 -283
rect 326 -322 328 -283
rect 338 -322 340 -283
rect 350 -322 352 -283
rect 375 -302 377 -282
rect 1330 -277 1332 -274
rect 1342 -277 1344 -274
rect 1365 -277 1367 -274
rect 1398 -277 1400 -274
rect 1430 -277 1432 -274
rect 965 -293 967 -288
rect 1093 -300 1095 -288
rect 1105 -307 1107 -288
rect 1117 -300 1119 -288
rect 1129 -307 1131 -288
rect 375 -317 377 -312
rect 314 -335 316 -332
rect 326 -335 328 -332
rect 338 -335 340 -332
rect 350 -335 352 -332
rect 1093 -333 1095 -325
rect 1105 -333 1107 -318
rect 1117 -333 1119 -326
rect 1129 -333 1131 -317
rect 1330 -318 1332 -297
rect 1330 -331 1332 -328
rect -305 -342 -303 -339
rect -293 -342 -291 -339
rect -281 -342 -279 -339
rect -269 -342 -267 -339
rect -601 -355 -599 -352
rect -589 -355 -587 -352
rect -566 -355 -564 -352
rect -533 -355 -531 -352
rect -501 -355 -499 -352
rect -601 -396 -599 -375
rect -601 -409 -599 -406
rect -589 -419 -587 -375
rect -566 -396 -564 -375
rect -554 -396 -552 -382
rect -533 -396 -531 -375
rect -521 -396 -519 -393
rect -501 -396 -499 -375
rect 27 -364 29 -339
rect 39 -364 41 -339
rect 64 -358 66 -338
rect 967 -354 969 -351
rect 1342 -341 1344 -297
rect 1365 -318 1367 -297
rect 1377 -318 1379 -304
rect 1398 -318 1400 -297
rect 1410 -318 1412 -315
rect 1430 -318 1432 -297
rect 1365 -341 1367 -328
rect 1377 -331 1379 -328
rect 1398 -331 1400 -328
rect 1410 -341 1412 -328
rect 1430 -331 1432 -328
rect 1342 -343 1412 -341
rect -305 -394 -303 -382
rect -293 -401 -291 -382
rect -281 -394 -279 -382
rect -269 -401 -267 -382
rect 64 -373 66 -368
rect 1093 -356 1095 -353
rect 1105 -356 1107 -353
rect 1117 -356 1119 -353
rect 1129 -356 1131 -353
rect 27 -388 29 -384
rect 39 -388 41 -384
rect 967 -394 969 -374
rect 170 -402 172 -398
rect 182 -402 184 -398
rect 207 -401 209 -398
rect -566 -419 -564 -406
rect -554 -409 -552 -406
rect -533 -409 -531 -406
rect -521 -419 -519 -406
rect -501 -409 -499 -406
rect -438 -409 -436 -406
rect -589 -421 -519 -419
rect -305 -427 -303 -419
rect -293 -427 -291 -412
rect -281 -427 -279 -420
rect -269 -427 -267 -411
rect 967 -409 969 -404
rect -438 -449 -436 -429
rect 170 -447 172 -422
rect 182 -447 184 -422
rect 207 -441 209 -421
rect -305 -450 -303 -447
rect -293 -450 -291 -447
rect -281 -450 -279 -447
rect -269 -450 -267 -447
rect -438 -464 -436 -459
rect 207 -456 209 -451
rect 170 -471 172 -467
rect 182 -471 184 -467
rect -435 -658 -433 -655
rect -435 -698 -433 -678
rect 138 -693 140 -690
rect 150 -693 152 -690
rect 162 -693 164 -690
rect -602 -714 -600 -711
rect -590 -714 -588 -711
rect -567 -714 -565 -711
rect -534 -714 -532 -711
rect -502 -714 -500 -711
rect -435 -713 -433 -708
rect -380 -727 -378 -723
rect -368 -727 -366 -723
rect -343 -726 -341 -723
rect -602 -755 -600 -734
rect -602 -768 -600 -765
rect -590 -778 -588 -734
rect -567 -755 -565 -734
rect -555 -755 -553 -741
rect -534 -755 -532 -734
rect -522 -755 -520 -752
rect -502 -755 -500 -734
rect -567 -778 -565 -765
rect -555 -768 -553 -765
rect -534 -768 -532 -765
rect -522 -778 -520 -765
rect -502 -768 -500 -765
rect -380 -772 -378 -747
rect -368 -772 -366 -747
rect -343 -766 -341 -746
rect -83 -756 -81 -752
rect -71 -756 -69 -752
rect -46 -755 -44 -752
rect 187 -729 189 -726
rect 927 -747 929 -744
rect -590 -780 -520 -778
rect -343 -781 -341 -776
rect -380 -796 -378 -792
rect -368 -796 -366 -792
rect -303 -803 -301 -800
rect -291 -803 -289 -800
rect -279 -803 -277 -800
rect -267 -803 -265 -800
rect -83 -801 -81 -776
rect -71 -801 -69 -776
rect -46 -795 -44 -775
rect 138 -789 140 -753
rect 150 -789 152 -753
rect 162 -789 164 -753
rect 187 -769 189 -749
rect 1055 -757 1057 -754
rect 1067 -757 1069 -754
rect 1079 -757 1081 -754
rect 1091 -757 1093 -754
rect 187 -784 189 -779
rect 927 -787 929 -767
rect -600 -817 -598 -814
rect -588 -817 -586 -814
rect -565 -817 -563 -814
rect -532 -817 -530 -814
rect -500 -817 -498 -814
rect -600 -858 -598 -837
rect -600 -871 -598 -868
rect -588 -881 -586 -837
rect -565 -858 -563 -837
rect -553 -858 -551 -844
rect -532 -858 -530 -837
rect -520 -858 -518 -855
rect -500 -858 -498 -837
rect 138 -802 140 -799
rect 150 -802 152 -799
rect 162 -802 164 -799
rect 927 -802 929 -797
rect -46 -810 -44 -805
rect 1055 -809 1057 -797
rect 1067 -816 1069 -797
rect 1079 -809 1081 -797
rect 1091 -816 1093 -797
rect 1333 -813 1335 -810
rect 1345 -813 1347 -810
rect 1368 -813 1370 -810
rect 1401 -813 1403 -810
rect 1433 -813 1435 -810
rect -83 -825 -81 -821
rect -71 -825 -69 -821
rect 1055 -842 1057 -834
rect 1067 -842 1069 -827
rect 1079 -842 1081 -835
rect 1091 -842 1093 -826
rect -303 -855 -301 -843
rect -291 -862 -289 -843
rect -279 -855 -277 -843
rect -267 -862 -265 -843
rect 18 -848 20 -844
rect 30 -848 32 -844
rect 55 -847 57 -844
rect -565 -881 -563 -868
rect -553 -871 -551 -868
rect -532 -871 -530 -868
rect -520 -881 -518 -868
rect -500 -871 -498 -868
rect -436 -870 -434 -867
rect 929 -863 931 -860
rect 1333 -854 1335 -833
rect -588 -883 -518 -881
rect -303 -888 -301 -880
rect -291 -888 -289 -873
rect -279 -888 -277 -881
rect -267 -888 -265 -872
rect -436 -910 -434 -890
rect 18 -893 20 -868
rect 30 -893 32 -868
rect 55 -887 57 -867
rect 1055 -865 1057 -862
rect 1067 -865 1069 -862
rect 1079 -865 1081 -862
rect 1091 -865 1093 -862
rect 1333 -867 1335 -864
rect 1345 -877 1347 -833
rect 1368 -854 1370 -833
rect 1380 -854 1382 -840
rect 1401 -854 1403 -833
rect 1413 -854 1415 -851
rect 1433 -854 1435 -833
rect 1368 -877 1370 -864
rect 1380 -867 1382 -864
rect 1401 -867 1403 -864
rect 1413 -877 1415 -864
rect 1433 -867 1435 -864
rect 1345 -879 1415 -877
rect -303 -911 -301 -908
rect -291 -911 -289 -908
rect -279 -911 -277 -908
rect -267 -911 -265 -908
rect 55 -902 57 -897
rect 929 -903 931 -883
rect 18 -917 20 -913
rect 30 -917 32 -913
rect 929 -918 931 -913
rect -436 -925 -434 -920
rect -682 -1021 -680 -1018
rect -670 -1021 -668 -1018
rect -647 -1021 -645 -1018
rect -614 -1021 -612 -1018
rect -582 -1021 -580 -1018
rect -682 -1062 -680 -1041
rect -682 -1075 -680 -1072
rect -670 -1085 -668 -1041
rect -647 -1062 -645 -1041
rect -635 -1062 -633 -1048
rect -614 -1062 -612 -1041
rect -602 -1062 -600 -1059
rect -582 -1062 -580 -1041
rect -647 -1085 -645 -1072
rect -635 -1075 -633 -1072
rect -614 -1075 -612 -1072
rect -602 -1085 -600 -1072
rect -582 -1075 -580 -1072
rect -670 -1087 -600 -1085
rect -434 -1112 -432 -1109
rect -434 -1152 -432 -1132
rect -600 -1164 -598 -1161
rect -588 -1164 -586 -1161
rect -565 -1164 -563 -1161
rect -532 -1164 -530 -1161
rect -500 -1164 -498 -1161
rect -434 -1167 -432 -1162
rect -110 -1163 -108 -1159
rect -98 -1163 -96 -1159
rect -73 -1162 -71 -1159
rect -379 -1181 -377 -1177
rect -367 -1181 -365 -1177
rect -342 -1180 -340 -1177
rect -600 -1205 -598 -1184
rect -600 -1218 -598 -1215
rect -588 -1228 -586 -1184
rect -565 -1205 -563 -1184
rect -553 -1205 -551 -1191
rect -532 -1205 -530 -1184
rect -520 -1205 -518 -1202
rect -500 -1205 -498 -1184
rect 903 -1170 905 -1167
rect -565 -1228 -563 -1215
rect -553 -1218 -551 -1215
rect -532 -1218 -530 -1215
rect -520 -1228 -518 -1215
rect -500 -1218 -498 -1215
rect -379 -1226 -377 -1201
rect -367 -1226 -365 -1201
rect -342 -1220 -340 -1200
rect -110 -1208 -108 -1183
rect -98 -1208 -96 -1183
rect -73 -1202 -71 -1182
rect 1031 -1180 1033 -1177
rect 1043 -1180 1045 -1177
rect 1055 -1180 1057 -1177
rect 1067 -1180 1069 -1177
rect -588 -1230 -518 -1228
rect 903 -1210 905 -1190
rect -73 -1217 -71 -1212
rect 903 -1225 905 -1220
rect -342 -1235 -340 -1230
rect -110 -1232 -108 -1228
rect -98 -1232 -96 -1228
rect 1031 -1232 1033 -1220
rect 6 -1240 8 -1237
rect 18 -1240 20 -1237
rect 1043 -1239 1045 -1220
rect 1055 -1232 1057 -1220
rect 1067 -1239 1069 -1220
rect 1325 -1223 1327 -1220
rect 1337 -1223 1339 -1220
rect 1360 -1223 1362 -1220
rect 1393 -1223 1395 -1220
rect 1425 -1223 1427 -1220
rect -379 -1250 -377 -1246
rect -367 -1250 -365 -1246
rect -302 -1257 -300 -1254
rect -290 -1257 -288 -1254
rect -278 -1257 -276 -1254
rect -266 -1257 -264 -1254
rect -599 -1274 -597 -1271
rect -587 -1274 -585 -1271
rect -564 -1274 -562 -1271
rect -531 -1274 -529 -1271
rect -499 -1274 -497 -1271
rect -599 -1315 -597 -1294
rect -599 -1328 -597 -1325
rect -587 -1338 -585 -1294
rect -564 -1315 -562 -1294
rect -552 -1315 -550 -1301
rect -531 -1315 -529 -1294
rect -519 -1315 -517 -1312
rect -499 -1315 -497 -1294
rect 43 -1258 45 -1255
rect 1031 -1265 1033 -1257
rect 1043 -1265 1045 -1250
rect 1055 -1265 1057 -1258
rect 1067 -1265 1069 -1249
rect 1325 -1264 1327 -1243
rect -302 -1309 -300 -1297
rect -290 -1316 -288 -1297
rect -278 -1309 -276 -1297
rect -266 -1316 -264 -1297
rect 6 -1304 8 -1280
rect 18 -1304 20 -1280
rect 43 -1298 45 -1278
rect 905 -1286 907 -1283
rect 1325 -1277 1327 -1274
rect 1031 -1288 1033 -1285
rect 1043 -1288 1045 -1285
rect 1055 -1288 1057 -1285
rect 1067 -1288 1069 -1285
rect 1337 -1287 1339 -1243
rect 1360 -1264 1362 -1243
rect 1372 -1264 1374 -1250
rect 1393 -1264 1395 -1243
rect 1405 -1264 1407 -1261
rect 1425 -1264 1427 -1243
rect 1360 -1287 1362 -1274
rect 1372 -1277 1374 -1274
rect 1393 -1277 1395 -1274
rect 1405 -1287 1407 -1274
rect 1425 -1277 1427 -1274
rect 1337 -1289 1407 -1287
rect 43 -1313 45 -1308
rect 6 -1317 8 -1314
rect 18 -1317 20 -1314
rect -435 -1324 -433 -1321
rect -564 -1338 -562 -1325
rect -552 -1328 -550 -1325
rect -531 -1328 -529 -1325
rect -519 -1338 -517 -1325
rect -499 -1328 -497 -1325
rect -587 -1340 -517 -1338
rect 905 -1326 907 -1306
rect -302 -1342 -300 -1334
rect -290 -1342 -288 -1327
rect -278 -1342 -276 -1335
rect -266 -1342 -264 -1326
rect 905 -1341 907 -1336
rect -435 -1364 -433 -1344
rect -302 -1365 -300 -1362
rect -290 -1365 -288 -1362
rect -278 -1365 -276 -1362
rect -266 -1365 -264 -1362
rect -435 -1379 -433 -1374
<< polycontact >>
rect 1335 932 1339 936
rect 1347 939 1351 943
rect 1382 938 1386 942
rect 1403 938 1407 942
rect 1435 938 1439 942
rect -440 615 -436 619
rect -602 556 -598 560
rect -590 563 -586 567
rect -555 562 -551 566
rect -534 562 -530 566
rect -502 562 -498 566
rect -139 573 -134 577
rect -386 549 -381 553
rect -375 540 -369 544
rect -348 547 -344 551
rect -128 564 -122 568
rect -101 571 -97 575
rect 970 585 974 589
rect 373 559 377 563
rect -604 454 -600 458
rect -592 461 -588 465
rect -557 460 -553 464
rect -536 460 -532 464
rect -504 460 -500 464
rect 392 550 396 554
rect 404 543 408 547
rect 416 536 420 540
rect 428 529 432 533
rect 440 522 444 526
rect 1098 559 1102 563
rect 465 538 469 542
rect 1110 552 1114 556
rect 1128 559 1132 563
rect 1140 552 1144 556
rect 1329 546 1333 550
rect 1341 553 1345 557
rect 1110 535 1114 539
rect 1098 528 1102 532
rect 1128 528 1132 532
rect 1140 535 1144 539
rect 1376 552 1380 556
rect 1397 552 1401 556
rect 1429 552 1433 556
rect -66 479 -61 483
rect -55 470 -49 474
rect -28 477 -24 481
rect -308 454 -304 458
rect -296 447 -292 451
rect -278 454 -274 458
rect -266 447 -262 451
rect 972 469 976 473
rect -296 430 -292 434
rect -308 423 -304 427
rect -278 423 -274 427
rect -266 430 -262 434
rect -441 403 -437 407
rect 20 378 25 382
rect 31 369 37 373
rect 58 376 62 380
rect 125 358 130 362
rect 136 349 142 353
rect 163 356 167 360
rect 251 299 256 303
rect 262 290 268 294
rect 289 297 293 301
rect -440 215 -436 219
rect -602 156 -598 160
rect -590 163 -586 167
rect -555 162 -551 166
rect -534 162 -530 166
rect -502 162 -498 166
rect -106 166 -101 170
rect -386 149 -381 153
rect -375 140 -369 144
rect -348 147 -344 151
rect -95 157 -89 161
rect -68 164 -64 168
rect 970 185 974 189
rect 364 148 368 152
rect -604 54 -600 58
rect -592 61 -588 65
rect -557 60 -553 64
rect -536 60 -532 64
rect -504 60 -500 64
rect 376 141 380 145
rect 388 134 392 138
rect 400 127 404 131
rect 412 120 416 124
rect 1098 159 1102 163
rect 1110 152 1114 156
rect 1128 159 1132 163
rect 1140 152 1144 156
rect 1329 146 1333 150
rect 1341 153 1345 157
rect 437 126 441 130
rect 1110 135 1114 139
rect 1098 128 1102 132
rect 1128 128 1132 132
rect 1140 135 1144 139
rect 1376 152 1380 156
rect 1397 152 1401 156
rect 1429 152 1433 156
rect 13 85 18 89
rect 24 76 30 80
rect 51 83 55 87
rect -308 54 -304 58
rect -296 47 -292 51
rect -278 54 -274 58
rect 972 69 976 73
rect -266 47 -262 51
rect -296 30 -292 34
rect -308 23 -304 27
rect -278 23 -274 27
rect -266 30 -262 34
rect -441 3 -437 7
rect 128 -11 133 -7
rect 139 -20 145 -16
rect 166 -13 170 -9
rect 256 -98 261 -94
rect 267 -107 273 -103
rect 294 -100 298 -96
rect -441 -232 -437 -228
rect -604 -291 -600 -287
rect -592 -284 -588 -280
rect -557 -285 -553 -281
rect -536 -285 -532 -281
rect -504 -285 -500 -281
rect -109 -279 -104 -275
rect -387 -298 -382 -294
rect -376 -307 -370 -303
rect -349 -300 -345 -296
rect -98 -288 -92 -284
rect -71 -281 -67 -277
rect 961 -273 965 -269
rect 309 -317 314 -313
rect 321 -310 326 -306
rect 333 -303 338 -299
rect 345 -296 350 -292
rect 371 -297 375 -293
rect 1089 -299 1093 -295
rect 1101 -306 1105 -302
rect 1119 -299 1123 -295
rect 1131 -306 1135 -302
rect 1326 -315 1330 -311
rect 1101 -323 1105 -319
rect 1089 -330 1093 -326
rect 1119 -330 1123 -326
rect 1338 -308 1342 -304
rect 1131 -323 1135 -319
rect -605 -393 -601 -389
rect -593 -386 -589 -382
rect -558 -387 -554 -383
rect -537 -387 -533 -383
rect -505 -387 -501 -383
rect 22 -351 27 -347
rect 33 -360 39 -356
rect 60 -353 64 -349
rect 1373 -309 1377 -305
rect 1394 -309 1398 -305
rect 1426 -309 1430 -305
rect -309 -393 -305 -389
rect -297 -400 -293 -396
rect -279 -393 -275 -389
rect 963 -389 967 -385
rect -267 -400 -263 -396
rect -297 -417 -293 -413
rect -309 -424 -305 -420
rect -279 -424 -275 -420
rect -267 -417 -263 -413
rect -442 -444 -438 -440
rect 165 -434 170 -430
rect 176 -443 182 -439
rect 203 -436 207 -432
rect -439 -693 -435 -689
rect -606 -752 -602 -748
rect -594 -745 -590 -741
rect -559 -746 -555 -742
rect -538 -746 -534 -742
rect -506 -746 -502 -742
rect -385 -759 -380 -755
rect -374 -768 -368 -764
rect -347 -761 -343 -757
rect 133 -765 138 -761
rect -88 -788 -83 -784
rect -77 -797 -71 -793
rect -50 -790 -46 -786
rect 145 -772 150 -768
rect 157 -779 162 -775
rect 183 -764 187 -760
rect 923 -782 927 -778
rect -604 -855 -600 -851
rect -592 -848 -588 -844
rect -557 -849 -553 -845
rect -536 -849 -532 -845
rect -504 -849 -500 -845
rect 1051 -808 1055 -804
rect 1063 -815 1067 -811
rect 1081 -808 1085 -804
rect 1093 -815 1097 -811
rect 1063 -832 1067 -828
rect 1051 -839 1055 -835
rect 1081 -839 1085 -835
rect 1093 -832 1097 -828
rect -307 -854 -303 -850
rect -295 -861 -291 -857
rect -277 -854 -273 -850
rect -265 -861 -261 -857
rect 1329 -851 1333 -847
rect 1341 -844 1345 -840
rect -295 -878 -291 -874
rect -307 -885 -303 -881
rect -277 -885 -273 -881
rect -265 -878 -261 -874
rect 13 -880 18 -876
rect -440 -905 -436 -901
rect 24 -889 30 -885
rect 51 -882 55 -878
rect 1376 -845 1380 -841
rect 1397 -845 1401 -841
rect 1429 -845 1433 -841
rect 925 -898 929 -894
rect -686 -1059 -682 -1055
rect -674 -1052 -670 -1048
rect -639 -1053 -635 -1049
rect -618 -1053 -614 -1049
rect -586 -1053 -582 -1049
rect -438 -1147 -434 -1143
rect -604 -1202 -600 -1198
rect -592 -1195 -588 -1191
rect -557 -1196 -553 -1192
rect -536 -1196 -532 -1192
rect -504 -1196 -500 -1192
rect -115 -1195 -110 -1191
rect -384 -1213 -379 -1209
rect -373 -1222 -367 -1218
rect -346 -1215 -342 -1211
rect -104 -1204 -98 -1200
rect -77 -1197 -73 -1193
rect 899 -1205 903 -1201
rect 1027 -1231 1031 -1227
rect 1039 -1238 1043 -1234
rect 1057 -1231 1061 -1227
rect 1069 -1238 1073 -1234
rect -603 -1312 -599 -1308
rect -591 -1305 -587 -1301
rect -556 -1306 -552 -1302
rect -535 -1306 -531 -1302
rect -503 -1306 -499 -1302
rect 1039 -1255 1043 -1251
rect 1027 -1262 1031 -1258
rect 1057 -1262 1061 -1258
rect 1069 -1255 1073 -1251
rect 1321 -1261 1325 -1257
rect 1333 -1254 1337 -1250
rect -306 -1308 -302 -1304
rect -294 -1315 -290 -1311
rect -276 -1308 -272 -1304
rect 1 -1301 6 -1297
rect 13 -1294 18 -1290
rect 39 -1293 43 -1289
rect -264 -1315 -260 -1311
rect 1368 -1255 1372 -1251
rect 1389 -1255 1393 -1251
rect 1421 -1255 1425 -1251
rect 901 -1321 905 -1317
rect -294 -1332 -290 -1328
rect -306 -1339 -302 -1335
rect -276 -1339 -272 -1335
rect -264 -1332 -260 -1328
rect -439 -1359 -435 -1355
<< metal1 >>
rect -638 1021 1527 1025
rect -638 567 -634 1021
rect 1319 943 1323 1021
rect 1338 974 1344 978
rect 1348 974 1354 978
rect 1358 974 1374 978
rect 1378 974 1402 978
rect 1406 974 1434 978
rect 1438 974 1452 978
rect 1334 970 1338 974
rect 1369 970 1373 974
rect 1402 970 1406 974
rect 1434 970 1438 974
rect 1381 950 1393 970
rect 1414 950 1426 970
rect 1319 939 1347 943
rect 1354 942 1358 950
rect 1389 942 1393 950
rect 1422 942 1426 950
rect 1442 942 1446 950
rect 1354 938 1382 942
rect 1389 938 1403 942
rect 1422 938 1435 942
rect 1442 938 1452 942
rect 1299 932 1335 936
rect 1299 930 1306 932
rect 1231 923 1306 930
rect 1354 929 1358 938
rect 1389 929 1393 938
rect 1422 929 1426 938
rect 1442 929 1446 938
rect 1346 919 1358 929
rect 1334 915 1338 919
rect 1369 915 1373 919
rect 1402 915 1406 919
rect 1434 915 1438 919
rect 1338 911 1369 915
rect 1373 911 1378 915
rect 1382 911 1389 915
rect 1393 911 1402 915
rect 1406 911 1412 915
rect 1416 911 1422 915
rect 1426 911 1434 915
rect 1438 911 1446 915
rect 372 709 468 710
rect 372 705 384 709
rect 392 705 400 709
rect 404 705 412 709
rect 416 705 424 709
rect 428 705 436 709
rect 440 705 446 709
rect 450 705 468 709
rect 372 704 468 705
rect 372 699 376 704
rect -448 656 -422 661
rect -441 650 -437 656
rect -433 619 -429 630
rect -475 615 -440 619
rect -433 615 -232 619
rect -599 598 -593 602
rect -589 598 -583 602
rect -579 598 -563 602
rect -559 598 -535 602
rect -531 598 -503 602
rect -499 598 -485 602
rect -603 594 -599 598
rect -568 594 -564 598
rect -535 594 -531 598
rect -503 594 -499 598
rect -556 574 -544 594
rect -523 574 -511 594
rect -638 563 -590 567
rect -583 566 -579 574
rect -548 566 -544 574
rect -515 566 -511 574
rect -495 566 -491 574
rect -475 566 -470 615
rect -433 610 -429 615
rect -441 594 -437 600
rect -441 590 -429 594
rect -386 592 -330 594
rect -638 465 -634 563
rect -583 562 -555 566
rect -548 562 -534 566
rect -515 562 -502 566
rect -495 562 -470 566
rect -609 556 -602 560
rect -583 553 -579 562
rect -548 553 -544 562
rect -515 553 -511 562
rect -495 553 -491 562
rect -591 543 -579 553
rect -475 556 -470 562
rect -386 588 -384 592
rect -380 588 -376 592
rect -372 588 -368 592
rect -364 588 -349 592
rect -345 588 -330 592
rect -386 586 -362 588
rect -386 581 -382 586
rect -366 581 -362 586
rect -349 582 -345 588
rect -475 549 -439 556
rect -432 553 -427 556
rect -378 554 -370 561
rect -432 549 -386 553
rect -378 551 -362 554
rect -341 551 -337 562
rect -378 550 -348 551
rect -366 547 -348 550
rect -341 547 -326 551
rect -603 539 -599 543
rect -568 539 -564 543
rect -535 539 -531 543
rect -503 539 -499 543
rect -474 540 -375 544
rect -599 535 -568 539
rect -564 535 -559 539
rect -555 535 -548 539
rect -544 535 -535 539
rect -531 535 -525 539
rect -521 535 -515 539
rect -511 535 -503 539
rect -499 535 -491 539
rect -601 496 -595 500
rect -591 496 -585 500
rect -581 496 -565 500
rect -561 496 -537 500
rect -533 496 -505 500
rect -501 496 -487 500
rect -605 492 -601 496
rect -570 492 -566 496
rect -537 492 -533 496
rect -505 492 -501 496
rect -558 472 -546 492
rect -525 472 -513 492
rect -638 461 -592 465
rect -585 464 -581 472
rect -550 464 -546 472
rect -517 464 -513 472
rect -497 464 -493 472
rect -474 488 -470 540
rect -366 536 -362 547
rect -341 542 -337 547
rect -349 526 -345 532
rect -386 511 -382 516
rect -349 511 -336 526
rect -392 507 -386 511
rect -382 507 -376 511
rect -372 507 -366 511
rect -362 507 -344 511
rect -340 507 -336 511
rect -326 521 -248 526
rect -326 488 -322 521
rect -474 484 -322 488
rect -305 510 -299 514
rect -295 510 -287 514
rect -283 510 -276 514
rect -272 510 -265 514
rect -309 509 -261 510
rect -309 505 -305 509
rect -265 505 -261 509
rect -474 464 -470 484
rect -638 167 -634 461
rect -585 460 -557 464
rect -550 460 -536 464
rect -517 460 -504 464
rect -497 460 -470 464
rect -611 454 -604 458
rect -585 451 -581 460
rect -550 451 -546 460
rect -517 451 -513 460
rect -497 451 -493 460
rect -593 441 -581 451
rect -605 437 -601 441
rect -570 437 -566 441
rect -537 437 -533 441
rect -505 437 -501 441
rect -601 433 -570 437
rect -566 433 -561 437
rect -557 433 -550 437
rect -546 433 -537 437
rect -533 433 -527 437
rect -523 433 -517 437
rect -513 433 -505 437
rect -501 433 -493 437
rect -475 407 -470 460
rect -432 455 -308 458
rect -449 444 -423 449
rect -442 438 -438 444
rect -340 434 -336 455
rect -320 454 -308 455
rect -308 447 -296 451
rect -289 443 -281 465
rect -252 458 -248 521
rect -274 454 -248 458
rect -236 454 -232 615
rect -139 616 -83 618
rect -139 612 -137 616
rect -133 612 -129 616
rect -125 612 -121 616
rect -117 612 -102 616
rect -98 612 -83 616
rect -139 610 -115 612
rect -139 605 -135 610
rect -119 605 -115 610
rect -102 606 -98 612
rect -131 578 -123 585
rect -195 573 -139 577
rect -131 575 -115 578
rect -94 575 -90 586
rect -131 574 -101 575
rect -195 570 -191 573
rect -262 447 -242 451
rect -234 447 -232 454
rect -210 566 -191 570
rect -119 571 -101 574
rect -94 571 327 575
rect -210 489 -206 566
rect -164 564 -128 568
rect -119 560 -115 571
rect -94 566 -90 571
rect -102 550 -98 556
rect 323 554 327 571
rect 341 563 345 631
rect 341 559 373 563
rect 323 550 392 554
rect -139 535 -135 540
rect -102 535 -89 550
rect 306 543 404 547
rect -145 531 -139 535
rect -135 531 -129 535
rect -125 531 -119 535
rect -115 531 -97 535
rect -93 531 -89 535
rect 29 539 310 543
rect -66 522 -10 524
rect -66 518 -64 522
rect -60 518 -56 522
rect -52 518 -48 522
rect -44 518 -29 522
rect -25 518 -10 522
rect -66 516 -42 518
rect -66 511 -62 516
rect -46 511 -42 516
rect -29 512 -25 518
rect -210 485 -84 489
rect -210 443 -206 485
rect -289 439 -205 443
rect -289 438 -213 439
rect -340 430 -296 434
rect -434 407 -430 418
rect -328 423 -308 427
rect -475 403 -441 407
rect -434 403 -363 407
rect -475 368 -470 403
rect -434 398 -430 403
rect -442 382 -438 388
rect -442 378 -430 382
rect -328 368 -323 423
rect -289 420 -281 438
rect -262 430 -242 434
rect -274 423 -252 427
rect -309 396 -305 400
rect -265 396 -261 400
rect -309 395 -261 396
rect -305 391 -299 395
rect -295 391 -287 395
rect -283 391 -275 395
rect -271 391 -265 395
rect -475 364 -323 368
rect -255 357 -252 423
rect -143 383 -139 485
rect -88 483 -84 485
rect -58 484 -50 491
rect -88 479 -66 483
rect -58 481 -42 484
rect -21 481 -17 492
rect 29 481 33 539
rect 313 536 416 540
rect 313 522 317 536
rect -58 480 -28 481
rect -46 477 -28 480
rect -21 477 33 481
rect 88 518 317 522
rect 321 529 428 533
rect 447 532 451 573
rect 464 586 468 704
rect 464 573 468 581
rect 472 542 476 553
rect 487 542 491 883
rect 852 695 860 698
rect 857 589 860 695
rect 938 641 1168 645
rect 938 589 942 641
rect 962 626 988 631
rect 969 620 973 626
rect 977 589 981 600
rect 1101 615 1107 619
rect 1111 615 1119 619
rect 1123 615 1130 619
rect 1134 615 1141 619
rect 1097 614 1145 615
rect 1097 610 1101 614
rect 1141 610 1145 614
rect 857 585 970 589
rect 977 585 1085 589
rect 977 580 981 585
rect 1059 582 1066 585
rect 969 564 973 570
rect 969 560 981 564
rect 1081 563 1085 585
rect 1081 559 1098 563
rect 455 538 465 542
rect 472 538 491 542
rect 1030 552 1110 556
rect 456 532 460 538
rect 472 533 476 538
rect 1030 536 1034 552
rect 1117 548 1125 570
rect 1164 563 1168 641
rect 1523 608 1527 1021
rect 1307 604 1527 608
rect 1132 559 1168 563
rect 1194 556 1199 559
rect 1144 552 1199 556
rect 1307 557 1311 604
rect 1332 588 1338 592
rect 1342 588 1348 592
rect 1352 588 1368 592
rect 1372 588 1396 592
rect 1400 588 1428 592
rect 1432 588 1446 592
rect 1328 584 1332 588
rect 1363 584 1367 588
rect 1396 584 1400 588
rect 1428 584 1432 588
rect 1375 564 1387 584
rect 1408 564 1420 584
rect 1307 553 1341 557
rect 1348 556 1352 564
rect 1383 556 1387 564
rect 1416 556 1420 564
rect 1436 556 1440 564
rect 1348 552 1376 556
rect 1383 552 1397 556
rect 1416 552 1429 556
rect 1436 552 1446 556
rect 1117 547 1219 548
rect 1314 547 1329 550
rect 1117 546 1329 547
rect 1117 543 1318 546
rect 1348 543 1352 552
rect 1383 543 1387 552
rect 1416 543 1420 552
rect 1436 543 1440 552
rect -117 470 -55 474
rect -352 348 -239 357
rect -117 305 -113 470
rect -46 466 -42 477
rect -21 472 -17 477
rect -29 456 -25 462
rect -66 441 -62 446
rect -29 441 -16 456
rect -72 437 -66 441
rect -62 437 -56 441
rect -52 437 -46 441
rect -42 437 -24 441
rect -20 437 -16 441
rect 20 421 76 423
rect 20 417 22 421
rect 26 417 30 421
rect 34 417 38 421
rect 42 417 57 421
rect 61 417 76 421
rect 20 415 44 417
rect 20 410 24 415
rect 40 410 44 415
rect 57 411 61 417
rect 28 383 36 390
rect 17 378 20 382
rect 28 380 44 383
rect 65 380 69 391
rect 88 380 92 518
rect 321 508 325 529
rect 447 528 460 532
rect 298 504 325 508
rect 329 522 440 526
rect 28 379 58 380
rect 40 376 58 379
rect 65 376 92 380
rect 125 401 181 403
rect 125 397 127 401
rect 131 397 135 401
rect 139 397 143 401
rect 147 397 162 401
rect 166 397 181 401
rect 125 395 149 397
rect 125 390 129 395
rect 145 390 149 395
rect -17 369 31 373
rect -117 301 -43 305
rect -448 256 -422 261
rect -441 250 -437 256
rect -433 219 -429 230
rect -475 215 -440 219
rect -433 215 -232 219
rect -599 198 -593 202
rect -589 198 -583 202
rect -579 198 -563 202
rect -559 198 -535 202
rect -531 198 -503 202
rect -499 198 -485 202
rect -603 194 -599 198
rect -568 194 -564 198
rect -535 194 -531 198
rect -503 194 -499 198
rect -556 174 -544 194
rect -523 174 -511 194
rect -638 163 -590 167
rect -583 166 -579 174
rect -548 166 -544 174
rect -515 166 -511 174
rect -495 166 -491 174
rect -475 166 -470 215
rect -433 210 -429 215
rect -441 194 -437 200
rect -441 190 -429 194
rect -386 192 -330 194
rect -638 65 -634 163
rect -583 162 -555 166
rect -548 162 -534 166
rect -515 162 -502 166
rect -495 162 -470 166
rect -609 156 -602 160
rect -583 153 -579 162
rect -548 153 -544 162
rect -515 153 -511 162
rect -495 153 -491 162
rect -591 143 -579 153
rect -475 156 -470 162
rect -386 188 -384 192
rect -380 188 -376 192
rect -372 188 -368 192
rect -364 188 -349 192
rect -345 188 -330 192
rect -386 186 -362 188
rect -386 181 -382 186
rect -366 181 -362 186
rect -349 182 -345 188
rect -475 149 -439 156
rect -432 153 -427 156
rect -378 154 -370 161
rect -432 149 -386 153
rect -378 151 -362 154
rect -341 151 -337 162
rect -378 150 -348 151
rect -366 147 -348 150
rect -341 147 -326 151
rect -603 139 -599 143
rect -568 139 -564 143
rect -535 139 -531 143
rect -503 139 -499 143
rect -474 140 -375 144
rect -599 135 -568 139
rect -564 135 -559 139
rect -555 135 -548 139
rect -544 135 -535 139
rect -531 135 -525 139
rect -521 135 -515 139
rect -511 135 -503 139
rect -499 135 -491 139
rect -601 96 -595 100
rect -591 96 -585 100
rect -581 96 -565 100
rect -561 96 -537 100
rect -533 96 -505 100
rect -501 96 -487 100
rect -605 92 -601 96
rect -570 92 -566 96
rect -537 92 -533 96
rect -505 92 -501 96
rect -558 72 -546 92
rect -525 72 -513 92
rect -638 61 -592 65
rect -585 64 -581 72
rect -550 64 -546 72
rect -517 64 -513 72
rect -497 64 -493 72
rect -474 88 -470 140
rect -366 136 -362 147
rect -341 142 -337 147
rect -349 126 -345 132
rect -386 111 -382 116
rect -349 111 -336 126
rect -392 107 -386 111
rect -382 107 -376 111
rect -372 107 -366 111
rect -362 107 -344 111
rect -340 107 -336 111
rect -326 121 -248 126
rect -326 88 -322 121
rect -474 84 -322 88
rect -305 110 -299 114
rect -295 110 -287 114
rect -283 110 -276 114
rect -272 110 -265 114
rect -309 109 -261 110
rect -309 105 -305 109
rect -265 105 -261 109
rect -474 64 -470 84
rect -638 -280 -634 61
rect -585 60 -557 64
rect -550 60 -536 64
rect -517 60 -504 64
rect -497 60 -470 64
rect -611 54 -604 58
rect -585 51 -581 60
rect -550 51 -546 60
rect -517 51 -513 60
rect -497 51 -493 60
rect -593 41 -581 51
rect -605 37 -601 41
rect -570 37 -566 41
rect -537 37 -533 41
rect -505 37 -501 41
rect -601 33 -570 37
rect -566 33 -561 37
rect -557 33 -550 37
rect -546 33 -537 37
rect -533 33 -527 37
rect -523 33 -517 37
rect -513 33 -505 37
rect -501 33 -493 37
rect -475 7 -470 60
rect -432 55 -308 58
rect -449 44 -423 49
rect -442 38 -438 44
rect -340 34 -336 55
rect -320 54 -308 55
rect -308 47 -296 51
rect -289 43 -281 65
rect -252 58 -248 121
rect -274 54 -248 58
rect -236 54 -232 215
rect -106 209 -50 211
rect -106 205 -104 209
rect -100 205 -96 209
rect -92 205 -88 209
rect -84 205 -69 209
rect -65 205 -50 209
rect -106 203 -82 205
rect -106 198 -102 203
rect -86 198 -82 203
rect -159 170 -155 183
rect -69 199 -65 205
rect -98 171 -90 178
rect -262 47 -242 51
rect -234 47 -232 54
rect -210 166 -106 170
rect -98 168 -82 171
rect -61 168 -57 179
rect -47 168 -43 301
rect -17 288 -13 369
rect 40 365 44 376
rect 65 371 69 376
rect 162 391 166 397
rect 133 363 141 370
rect 57 355 61 361
rect 120 358 125 362
rect 133 360 149 363
rect 170 360 174 371
rect 298 360 302 504
rect 329 500 333 522
rect 447 519 451 528
rect 372 514 451 519
rect 372 511 376 514
rect 399 511 407 514
rect 423 511 431 514
rect 447 511 451 514
rect 940 532 1034 536
rect 1066 535 1110 539
rect 464 515 468 523
rect 464 507 468 511
rect 455 502 468 507
rect 133 359 163 360
rect 145 356 163 359
rect 170 356 302 360
rect 321 496 333 500
rect 382 497 395 501
rect 411 497 419 501
rect 435 497 443 501
rect 457 497 462 502
rect 20 340 24 345
rect 57 340 70 355
rect 14 336 20 340
rect 24 336 30 340
rect 34 336 40 340
rect 44 336 62 340
rect 66 336 70 340
rect 98 349 136 353
rect -17 284 87 288
rect -98 167 -68 168
rect -210 89 -206 166
rect -86 164 -68 167
rect -61 164 58 168
rect 65 164 66 168
rect -179 157 -95 161
rect -179 155 -168 157
rect -86 153 -82 164
rect -61 159 -57 164
rect -69 143 -65 149
rect -106 128 -102 133
rect -69 128 -56 143
rect -112 124 -106 128
rect -102 124 -96 128
rect -92 124 -86 128
rect -82 124 -64 128
rect -60 124 -56 128
rect 13 128 69 130
rect 13 124 15 128
rect 19 124 23 128
rect 27 124 31 128
rect 35 124 50 128
rect 54 124 69 128
rect 13 122 37 124
rect 13 117 17 122
rect 33 117 37 122
rect 50 118 54 124
rect 21 90 29 97
rect -210 85 13 89
rect 21 87 37 90
rect 58 87 62 98
rect 83 87 87 284
rect 98 254 102 349
rect 145 345 149 356
rect 170 351 174 356
rect 251 342 307 344
rect 162 335 166 341
rect 251 338 253 342
rect 257 338 261 342
rect 265 338 269 342
rect 273 338 288 342
rect 292 338 307 342
rect 251 336 275 338
rect 125 320 129 325
rect 162 320 175 335
rect 119 316 125 320
rect 129 316 135 320
rect 139 316 145 320
rect 149 316 167 320
rect 171 316 175 320
rect 251 331 255 336
rect 271 331 275 336
rect 288 332 292 338
rect 259 304 267 311
rect 246 299 251 303
rect 259 301 275 304
rect 296 301 300 312
rect 321 301 325 496
rect 382 493 385 497
rect 391 496 462 497
rect 391 493 401 496
rect 382 492 401 493
rect 405 492 413 496
rect 417 492 425 496
rect 429 492 437 496
rect 441 492 447 496
rect 451 492 462 496
rect 940 473 944 532
rect 1082 528 1098 532
rect 964 510 990 515
rect 971 504 975 510
rect 979 473 983 484
rect 1082 473 1086 528
rect 1117 525 1125 543
rect 1144 535 1174 539
rect 1340 533 1352 543
rect 1132 528 1163 532
rect 1097 501 1101 505
rect 1141 501 1145 505
rect 1097 500 1145 501
rect 1101 496 1107 500
rect 1111 496 1119 500
rect 1123 496 1131 500
rect 1135 496 1141 500
rect 891 469 972 473
rect 979 469 1078 473
rect 891 461 895 469
rect 768 457 895 461
rect 940 432 944 469
rect 979 464 983 469
rect 971 448 975 454
rect 971 444 983 448
rect 1159 432 1163 528
rect 1328 529 1332 533
rect 1363 529 1367 533
rect 1396 529 1400 533
rect 1428 529 1432 533
rect 1332 525 1363 529
rect 1367 525 1372 529
rect 1376 525 1383 529
rect 1387 525 1396 529
rect 1400 525 1406 529
rect 1410 525 1416 529
rect 1420 525 1428 529
rect 1432 525 1440 529
rect 940 428 1163 432
rect 259 300 289 301
rect 271 297 289 300
rect 296 297 325 301
rect 204 290 262 294
rect 98 250 191 254
rect 128 164 161 168
rect 21 86 51 87
rect -210 43 -206 85
rect -289 39 -205 43
rect -289 38 -213 39
rect -340 30 -296 34
rect -434 7 -430 18
rect -328 23 -308 27
rect -475 3 -441 7
rect -434 3 -363 7
rect -475 -32 -470 3
rect -434 -2 -430 3
rect -442 -18 -438 -12
rect -442 -22 -430 -18
rect -328 -32 -323 23
rect -289 20 -281 38
rect -262 30 -242 34
rect -274 23 -252 27
rect -309 -4 -305 0
rect -265 -4 -261 0
rect -309 -5 -261 -4
rect -305 -9 -299 -5
rect -295 -9 -287 -5
rect -283 -9 -275 -5
rect -271 -9 -265 -5
rect -475 -36 -323 -32
rect -255 -43 -252 23
rect -102 14 -95 85
rect 33 83 51 86
rect 58 83 163 87
rect -46 76 24 80
rect -352 -52 -239 -43
rect -449 -191 -423 -186
rect -442 -197 -438 -191
rect -434 -228 -430 -217
rect -476 -232 -441 -228
rect -434 -232 -233 -228
rect -601 -249 -595 -245
rect -591 -249 -585 -245
rect -581 -249 -565 -245
rect -561 -249 -537 -245
rect -533 -249 -505 -245
rect -501 -249 -487 -245
rect -605 -253 -601 -249
rect -570 -253 -566 -249
rect -537 -253 -533 -249
rect -505 -253 -501 -249
rect -558 -273 -546 -253
rect -525 -273 -513 -253
rect -638 -284 -592 -280
rect -585 -281 -581 -273
rect -550 -281 -546 -273
rect -517 -281 -513 -273
rect -497 -281 -493 -273
rect -476 -281 -471 -232
rect -434 -237 -430 -232
rect -442 -253 -438 -247
rect -442 -257 -430 -253
rect -387 -255 -331 -253
rect -638 -382 -634 -284
rect -585 -285 -557 -281
rect -550 -285 -536 -281
rect -517 -285 -504 -281
rect -497 -285 -471 -281
rect -611 -291 -604 -287
rect -585 -294 -581 -285
rect -550 -294 -546 -285
rect -517 -294 -513 -285
rect -497 -294 -493 -285
rect -593 -304 -581 -294
rect -476 -291 -471 -285
rect -387 -259 -385 -255
rect -381 -259 -377 -255
rect -373 -259 -369 -255
rect -365 -259 -350 -255
rect -346 -259 -331 -255
rect -387 -261 -363 -259
rect -387 -266 -383 -261
rect -367 -266 -363 -261
rect -350 -265 -346 -259
rect -476 -298 -440 -291
rect -433 -294 -428 -291
rect -379 -293 -371 -286
rect -433 -298 -387 -294
rect -379 -296 -363 -293
rect -342 -296 -338 -285
rect -379 -297 -349 -296
rect -367 -300 -349 -297
rect -342 -300 -312 -296
rect -605 -308 -601 -304
rect -570 -308 -566 -304
rect -537 -308 -533 -304
rect -505 -308 -501 -304
rect -475 -307 -376 -303
rect -601 -312 -570 -308
rect -566 -312 -561 -308
rect -557 -312 -550 -308
rect -546 -312 -537 -308
rect -533 -312 -527 -308
rect -523 -312 -517 -308
rect -513 -312 -505 -308
rect -501 -312 -493 -308
rect -602 -351 -596 -347
rect -592 -351 -586 -347
rect -582 -351 -566 -347
rect -562 -351 -538 -347
rect -534 -351 -506 -347
rect -502 -351 -488 -347
rect -606 -355 -602 -351
rect -571 -355 -567 -351
rect -538 -355 -534 -351
rect -506 -355 -502 -351
rect -559 -375 -547 -355
rect -526 -375 -514 -355
rect -638 -386 -593 -382
rect -586 -383 -582 -375
rect -551 -383 -547 -375
rect -518 -383 -514 -375
rect -498 -383 -494 -375
rect -475 -359 -471 -307
rect -367 -311 -363 -300
rect -342 -305 -338 -300
rect -350 -321 -346 -315
rect -387 -336 -383 -331
rect -350 -336 -337 -321
rect -393 -340 -387 -336
rect -383 -340 -377 -336
rect -373 -340 -367 -336
rect -363 -340 -345 -336
rect -341 -340 -337 -336
rect -327 -326 -249 -321
rect -327 -359 -323 -326
rect -475 -363 -323 -359
rect -306 -337 -300 -333
rect -296 -337 -288 -333
rect -284 -337 -277 -333
rect -273 -337 -266 -333
rect -310 -338 -262 -337
rect -310 -342 -306 -338
rect -266 -342 -262 -338
rect -475 -383 -471 -363
rect -638 -741 -634 -386
rect -586 -387 -558 -383
rect -551 -387 -537 -383
rect -518 -387 -505 -383
rect -498 -387 -471 -383
rect -612 -393 -605 -389
rect -586 -396 -582 -387
rect -551 -396 -547 -387
rect -518 -396 -514 -387
rect -498 -396 -494 -387
rect -594 -406 -582 -396
rect -606 -410 -602 -406
rect -571 -410 -567 -406
rect -538 -410 -534 -406
rect -506 -410 -502 -406
rect -602 -414 -571 -410
rect -567 -414 -562 -410
rect -558 -414 -551 -410
rect -547 -414 -538 -410
rect -534 -414 -528 -410
rect -524 -414 -518 -410
rect -514 -414 -506 -410
rect -502 -414 -494 -410
rect -476 -440 -471 -387
rect -433 -392 -309 -389
rect -450 -403 -424 -398
rect -443 -409 -439 -403
rect -341 -413 -337 -392
rect -321 -393 -309 -392
rect -309 -400 -297 -396
rect -290 -404 -282 -382
rect -253 -389 -249 -326
rect -275 -393 -249 -389
rect -237 -393 -233 -232
rect -109 -236 -53 -234
rect -109 -240 -107 -236
rect -103 -240 -99 -236
rect -95 -240 -91 -236
rect -87 -240 -72 -236
rect -68 -240 -53 -236
rect -109 -242 -85 -240
rect -109 -247 -105 -242
rect -89 -247 -85 -242
rect -72 -246 -68 -240
rect -101 -274 -93 -267
rect -263 -400 -243 -396
rect -235 -400 -233 -393
rect -187 -279 -109 -275
rect -101 -277 -85 -274
rect -64 -277 -60 -266
rect -46 -277 -42 76
rect 33 72 37 83
rect 58 78 62 83
rect 50 62 54 68
rect 13 47 17 52
rect 50 47 63 62
rect 7 43 13 47
rect 17 43 23 47
rect 27 43 33 47
rect 37 43 55 47
rect 59 43 63 47
rect 128 32 184 34
rect 128 28 130 32
rect 134 28 138 32
rect 142 28 146 32
rect 150 28 165 32
rect 169 28 184 32
rect 128 26 152 28
rect 128 21 132 26
rect 148 21 152 26
rect 98 0 105 7
rect 165 22 169 28
rect 100 -7 105 0
rect 136 -6 144 1
rect 100 -11 128 -7
rect 136 -9 152 -6
rect 173 -9 177 2
rect 187 -9 191 250
rect 204 28 208 290
rect 271 286 275 297
rect 296 292 300 297
rect 288 276 292 282
rect 251 261 255 266
rect 288 261 301 276
rect 245 257 251 261
rect 255 257 261 261
rect 265 257 271 261
rect 275 257 293 261
rect 297 257 301 261
rect 363 270 440 271
rect 367 266 372 270
rect 376 266 384 270
rect 388 266 396 270
rect 400 266 408 270
rect 412 266 418 270
rect 422 266 440 270
rect 363 265 440 266
rect 363 261 367 265
rect 313 218 318 223
rect 237 164 292 168
rect 288 145 292 164
rect 314 152 318 218
rect 314 148 364 152
rect 288 141 376 145
rect 267 134 388 138
rect 267 87 271 134
rect 238 83 271 87
rect 296 127 400 131
rect 419 130 423 161
rect 436 174 440 265
rect 938 241 1168 245
rect 886 185 888 189
rect 938 189 942 241
rect 962 226 988 231
rect 969 220 973 226
rect 977 189 981 200
rect 1101 215 1107 219
rect 1111 215 1119 219
rect 1123 215 1130 219
rect 1134 215 1141 219
rect 1097 214 1145 215
rect 1097 210 1101 214
rect 1141 210 1145 214
rect 894 185 970 189
rect 977 185 1085 189
rect 977 180 981 185
rect 436 161 440 169
rect 1059 182 1066 185
rect 969 164 973 170
rect 969 160 981 164
rect 1081 163 1085 185
rect 1081 159 1098 163
rect 444 130 448 141
rect 1030 152 1110 156
rect 1030 136 1034 152
rect 1117 148 1125 170
rect 1164 163 1168 241
rect 1523 208 1527 604
rect 1307 204 1527 208
rect 1132 159 1168 163
rect 1194 156 1199 159
rect 1144 152 1199 156
rect 1307 157 1311 204
rect 1332 188 1338 192
rect 1342 188 1348 192
rect 1352 188 1368 192
rect 1372 188 1396 192
rect 1400 188 1428 192
rect 1432 188 1446 192
rect 1328 184 1332 188
rect 1363 184 1367 188
rect 1396 184 1400 188
rect 1428 184 1432 188
rect 1375 164 1387 184
rect 1408 164 1420 184
rect 1307 153 1341 157
rect 1348 156 1352 164
rect 1383 156 1387 164
rect 1416 156 1420 164
rect 1436 156 1440 164
rect 1348 152 1376 156
rect 1383 152 1397 156
rect 1416 152 1429 156
rect 1436 152 1446 156
rect 1117 147 1219 148
rect 1314 147 1329 150
rect 1117 146 1329 147
rect 1117 143 1318 146
rect 1348 143 1352 152
rect 1383 143 1387 152
rect 1416 143 1420 152
rect 1436 143 1440 152
rect 296 28 300 127
rect 419 126 437 130
rect 444 126 468 130
rect 940 132 1034 136
rect 1066 135 1110 139
rect 321 120 412 124
rect 321 28 325 120
rect 419 117 423 126
rect 444 121 448 126
rect 371 112 423 117
rect 371 109 379 112
rect 395 109 403 112
rect 419 109 423 112
rect 436 103 440 111
rect 363 95 367 99
rect 383 95 391 99
rect 407 95 415 99
rect 436 95 440 99
rect 363 94 440 95
rect 367 90 373 94
rect 377 90 385 94
rect 389 90 397 94
rect 401 90 409 94
rect 413 90 419 94
rect 423 90 440 94
rect 940 73 944 132
rect 1082 128 1098 132
rect 964 110 990 115
rect 971 104 975 110
rect 979 73 983 84
rect 1082 73 1086 128
rect 1117 125 1125 143
rect 1144 135 1174 139
rect 1340 133 1352 143
rect 1132 128 1163 132
rect 1097 101 1101 105
rect 1141 101 1145 105
rect 1097 100 1145 101
rect 1101 96 1107 100
rect 1111 96 1119 100
rect 1123 96 1131 100
rect 1135 96 1141 100
rect 891 69 972 73
rect 979 69 1078 73
rect 891 61 895 69
rect 204 24 325 28
rect 296 -9 300 24
rect 136 -10 166 -9
rect 148 -13 166 -10
rect 173 -13 300 -9
rect 84 -20 139 -16
rect 84 -277 88 -20
rect 148 -24 152 -13
rect 173 -18 177 -13
rect 165 -34 169 -28
rect 128 -49 132 -44
rect 165 -49 178 -34
rect 122 -53 128 -49
rect 132 -53 138 -49
rect 142 -53 148 -49
rect 152 -53 170 -49
rect 174 -53 178 -49
rect 256 -55 312 -53
rect 256 -59 258 -55
rect 262 -59 266 -55
rect 270 -59 274 -55
rect 278 -59 293 -55
rect 297 -59 312 -55
rect 256 -61 280 -59
rect 256 -66 260 -61
rect 276 -66 280 -61
rect 293 -65 297 -59
rect 264 -93 272 -86
rect 186 -98 256 -94
rect 264 -96 280 -93
rect 301 -96 305 -85
rect 321 -96 325 24
rect 264 -97 294 -96
rect 276 -100 294 -97
rect 301 -100 325 -96
rect 583 57 895 61
rect 228 -107 267 -103
rect 228 -246 235 -107
rect 276 -111 280 -100
rect 301 -105 305 -100
rect 293 -121 297 -115
rect 256 -136 260 -131
rect 293 -136 306 -121
rect 250 -140 256 -136
rect 260 -140 266 -136
rect 270 -140 276 -136
rect 280 -140 298 -136
rect 302 -140 306 -136
rect 313 -199 318 -195
rect 322 -199 330 -195
rect 334 -199 343 -195
rect 347 -199 353 -195
rect 357 -199 374 -195
rect 309 -203 313 -199
rect 261 -214 270 -212
rect 261 -218 293 -214
rect -101 -278 -71 -277
rect -187 -347 -182 -279
rect -89 -281 -71 -278
rect -64 -281 285 -277
rect -151 -288 -98 -284
rect -151 -290 -145 -288
rect -89 -292 -85 -281
rect -64 -286 -60 -281
rect -72 -302 -68 -296
rect -109 -317 -105 -312
rect -72 -317 -59 -302
rect -115 -321 -109 -317
rect -105 -321 -99 -317
rect -95 -321 -89 -317
rect -85 -321 -67 -317
rect -63 -321 -59 -317
rect 22 -308 78 -306
rect 22 -312 24 -308
rect 28 -312 32 -308
rect 36 -312 40 -308
rect 44 -312 59 -308
rect 63 -312 78 -308
rect 22 -314 46 -312
rect 22 -319 26 -314
rect 42 -319 46 -314
rect 59 -318 63 -312
rect 30 -346 38 -339
rect -187 -351 22 -347
rect 30 -349 46 -346
rect 67 -349 71 -338
rect 84 -349 88 -281
rect 281 -299 285 -281
rect 289 -292 293 -218
rect 370 -252 374 -199
rect 374 -256 388 -252
rect 370 -262 374 -256
rect 289 -296 345 -292
rect 353 -293 357 -283
rect 378 -293 382 -282
rect 583 -293 587 57
rect 940 32 944 69
rect 979 64 983 69
rect 971 48 975 54
rect 971 44 983 48
rect 1159 32 1163 128
rect 1328 129 1332 133
rect 1363 129 1367 133
rect 1396 129 1400 133
rect 1428 129 1432 133
rect 1332 125 1363 129
rect 1367 125 1372 129
rect 1376 125 1383 129
rect 1387 125 1396 129
rect 1400 125 1406 129
rect 1410 125 1416 129
rect 1420 125 1428 129
rect 1432 125 1440 129
rect 940 28 1163 32
rect 929 -217 1159 -213
rect 929 -269 933 -217
rect 953 -232 979 -227
rect 960 -238 964 -232
rect 968 -269 972 -258
rect 1092 -243 1098 -239
rect 1102 -243 1110 -239
rect 1114 -243 1121 -239
rect 1125 -243 1132 -239
rect 1088 -244 1136 -243
rect 1088 -248 1092 -244
rect 1132 -248 1136 -244
rect 887 -273 961 -269
rect 968 -273 1076 -269
rect 887 -274 916 -273
rect 887 -277 892 -274
rect 353 -297 371 -293
rect 378 -297 587 -293
rect 661 -282 892 -277
rect 968 -278 972 -273
rect 281 -303 333 -299
rect 195 -310 321 -306
rect 195 -349 199 -310
rect 353 -313 357 -297
rect 378 -302 382 -297
rect 30 -350 60 -349
rect -187 -404 -182 -351
rect -57 -355 -51 -351
rect 42 -353 60 -350
rect 67 -353 199 -349
rect 289 -317 309 -313
rect -27 -360 33 -356
rect -290 -409 -182 -404
rect -341 -417 -297 -413
rect -435 -440 -431 -429
rect -329 -424 -309 -420
rect -476 -444 -442 -440
rect -435 -444 -364 -440
rect -476 -479 -471 -444
rect -435 -449 -431 -444
rect -443 -465 -439 -459
rect -443 -469 -431 -465
rect -329 -479 -324 -424
rect -290 -427 -282 -409
rect -263 -417 -243 -413
rect -275 -424 -253 -420
rect -310 -451 -306 -447
rect -266 -451 -262 -447
rect -310 -452 -262 -451
rect -306 -456 -300 -452
rect -296 -456 -288 -452
rect -284 -456 -276 -452
rect -272 -456 -266 -452
rect -476 -483 -324 -479
rect -256 -490 -253 -424
rect -353 -499 -240 -490
rect -447 -652 -421 -647
rect -440 -658 -436 -652
rect -432 -689 -428 -678
rect -474 -693 -439 -689
rect -432 -693 -231 -689
rect -603 -710 -597 -706
rect -593 -710 -587 -706
rect -583 -710 -567 -706
rect -563 -710 -539 -706
rect -535 -710 -507 -706
rect -503 -710 -489 -706
rect -607 -714 -603 -710
rect -572 -714 -568 -710
rect -539 -714 -535 -710
rect -507 -714 -503 -710
rect -560 -734 -548 -714
rect -527 -734 -515 -714
rect -638 -745 -594 -741
rect -587 -742 -583 -734
rect -552 -742 -548 -734
rect -519 -742 -515 -734
rect -499 -742 -495 -734
rect -474 -742 -469 -693
rect -432 -698 -428 -693
rect -440 -714 -436 -708
rect -440 -718 -428 -714
rect -385 -716 -329 -714
rect -638 -844 -634 -745
rect -587 -746 -559 -742
rect -552 -746 -538 -742
rect -519 -746 -506 -742
rect -499 -746 -469 -742
rect -613 -752 -606 -748
rect -587 -755 -583 -746
rect -552 -755 -548 -746
rect -519 -755 -515 -746
rect -499 -755 -495 -746
rect -595 -765 -583 -755
rect -474 -752 -469 -746
rect -385 -720 -383 -716
rect -379 -720 -375 -716
rect -371 -720 -367 -716
rect -363 -720 -348 -716
rect -344 -720 -329 -716
rect -385 -722 -361 -720
rect -385 -727 -381 -722
rect -365 -727 -361 -722
rect -348 -726 -344 -720
rect -474 -759 -438 -752
rect -431 -755 -426 -752
rect -377 -754 -369 -747
rect -431 -759 -385 -755
rect -377 -757 -361 -754
rect -340 -757 -336 -746
rect -377 -758 -347 -757
rect -365 -761 -347 -758
rect -340 -761 -317 -757
rect -607 -769 -603 -765
rect -572 -769 -568 -765
rect -539 -769 -535 -765
rect -507 -769 -503 -765
rect -473 -768 -374 -764
rect -603 -773 -572 -769
rect -568 -773 -563 -769
rect -559 -773 -552 -769
rect -548 -773 -539 -769
rect -535 -773 -529 -769
rect -525 -773 -519 -769
rect -515 -773 -507 -769
rect -503 -773 -495 -769
rect -601 -813 -595 -809
rect -591 -813 -585 -809
rect -581 -813 -565 -809
rect -561 -813 -537 -809
rect -533 -813 -505 -809
rect -501 -813 -487 -809
rect -605 -817 -601 -813
rect -570 -817 -566 -813
rect -537 -817 -533 -813
rect -505 -817 -501 -813
rect -558 -837 -546 -817
rect -525 -837 -513 -817
rect -638 -848 -592 -844
rect -585 -845 -581 -837
rect -550 -845 -546 -837
rect -517 -845 -513 -837
rect -497 -845 -493 -837
rect -473 -820 -469 -768
rect -365 -772 -361 -761
rect -340 -766 -336 -761
rect -348 -782 -344 -776
rect -385 -797 -381 -792
rect -348 -797 -335 -782
rect -391 -801 -385 -797
rect -381 -801 -375 -797
rect -371 -801 -365 -797
rect -361 -801 -343 -797
rect -339 -801 -335 -797
rect -325 -787 -247 -782
rect -325 -820 -321 -787
rect -473 -824 -321 -820
rect -304 -798 -298 -794
rect -294 -798 -286 -794
rect -282 -798 -275 -794
rect -271 -798 -264 -794
rect -308 -799 -260 -798
rect -308 -803 -304 -799
rect -264 -803 -260 -799
rect -473 -845 -469 -824
rect -638 -980 -634 -848
rect -585 -849 -557 -845
rect -550 -849 -536 -845
rect -517 -849 -504 -845
rect -497 -849 -469 -845
rect -611 -855 -604 -851
rect -585 -858 -581 -849
rect -550 -858 -546 -849
rect -517 -858 -513 -849
rect -497 -858 -493 -849
rect -593 -868 -581 -858
rect -605 -872 -601 -868
rect -570 -872 -566 -868
rect -537 -872 -533 -868
rect -505 -872 -501 -868
rect -601 -876 -570 -872
rect -566 -876 -561 -872
rect -557 -876 -550 -872
rect -546 -876 -537 -872
rect -533 -876 -527 -872
rect -523 -876 -517 -872
rect -513 -876 -505 -872
rect -501 -876 -493 -872
rect -474 -901 -469 -849
rect -431 -853 -307 -850
rect -448 -864 -422 -859
rect -441 -870 -437 -864
rect -339 -874 -335 -853
rect -319 -854 -307 -853
rect -307 -861 -295 -857
rect -288 -865 -280 -843
rect -251 -850 -247 -787
rect -273 -854 -247 -850
rect -235 -854 -231 -693
rect -88 -745 -32 -743
rect -88 -749 -86 -745
rect -82 -749 -78 -745
rect -74 -749 -70 -745
rect -66 -749 -51 -745
rect -47 -749 -32 -745
rect -88 -751 -64 -749
rect -88 -756 -84 -751
rect -68 -756 -64 -751
rect -51 -755 -47 -749
rect -80 -783 -72 -776
rect -261 -861 -241 -857
rect -233 -861 -231 -854
rect -171 -788 -88 -784
rect -80 -786 -64 -783
rect -43 -786 -39 -775
rect -27 -786 -23 -360
rect 42 -364 46 -353
rect 67 -358 71 -353
rect 59 -374 63 -368
rect 22 -389 26 -384
rect 59 -389 72 -374
rect 16 -393 22 -389
rect 26 -393 32 -389
rect 36 -393 42 -389
rect 46 -393 64 -389
rect 68 -393 72 -389
rect 165 -391 221 -389
rect 165 -395 167 -391
rect 171 -395 175 -391
rect 179 -395 183 -391
rect 187 -395 202 -391
rect 206 -395 221 -391
rect 165 -397 189 -395
rect 165 -402 169 -397
rect 185 -402 189 -397
rect 202 -401 206 -395
rect 67 -430 74 -428
rect 173 -429 181 -422
rect 67 -434 165 -430
rect 173 -432 189 -429
rect 210 -432 214 -421
rect 289 -432 293 -317
rect 317 -319 357 -313
rect 317 -322 325 -319
rect 341 -322 349 -319
rect 370 -322 374 -312
rect 309 -336 313 -332
rect 329 -336 337 -332
rect 353 -336 357 -332
rect 370 -336 374 -326
rect 313 -340 319 -336
rect 323 -340 331 -336
rect 335 -340 343 -336
rect 347 -340 353 -336
rect 357 -340 374 -336
rect 173 -433 203 -432
rect 81 -533 86 -434
rect 185 -436 203 -433
rect 210 -436 293 -432
rect 115 -443 176 -439
rect 115 -446 135 -443
rect 185 -447 189 -436
rect 210 -441 214 -436
rect 202 -457 206 -451
rect 165 -472 169 -467
rect 202 -472 215 -457
rect 159 -476 165 -472
rect 169 -476 175 -472
rect 179 -476 185 -472
rect 189 -476 207 -472
rect 211 -476 215 -472
rect 661 -533 666 -282
rect 1050 -276 1057 -273
rect 960 -294 964 -288
rect 960 -298 972 -294
rect 1072 -295 1076 -273
rect 1072 -299 1089 -295
rect 1021 -306 1101 -302
rect 1021 -322 1025 -306
rect 1108 -310 1116 -288
rect 1155 -295 1159 -217
rect 1523 -252 1527 204
rect 1299 -256 1527 -252
rect 1123 -299 1159 -295
rect 1185 -302 1190 -299
rect 1135 -306 1190 -302
rect 1299 -304 1303 -256
rect 1329 -273 1335 -269
rect 1339 -273 1345 -269
rect 1349 -273 1365 -269
rect 1369 -273 1393 -269
rect 1397 -273 1425 -269
rect 1429 -273 1443 -269
rect 1325 -277 1329 -273
rect 1360 -277 1364 -273
rect 1393 -277 1397 -273
rect 1425 -277 1429 -273
rect 1372 -297 1384 -277
rect 1405 -297 1417 -277
rect 1299 -308 1338 -304
rect 1345 -305 1349 -297
rect 1380 -305 1384 -297
rect 1413 -305 1417 -297
rect 1433 -305 1437 -297
rect 1345 -309 1373 -305
rect 1380 -309 1394 -305
rect 1413 -309 1426 -305
rect 1433 -309 1443 -305
rect 1108 -311 1225 -310
rect 1108 -315 1326 -311
rect 931 -326 1025 -322
rect 1057 -323 1101 -319
rect 81 -538 666 -533
rect 780 -385 784 -382
rect 931 -385 935 -326
rect 1073 -330 1089 -326
rect 955 -348 981 -343
rect 962 -354 966 -348
rect 970 -385 974 -374
rect 1073 -385 1077 -330
rect 1108 -333 1116 -315
rect 1345 -318 1349 -309
rect 1380 -318 1384 -309
rect 1413 -318 1417 -309
rect 1433 -318 1437 -309
rect 1135 -323 1165 -319
rect 1123 -330 1154 -326
rect 1088 -357 1092 -353
rect 1132 -357 1136 -353
rect 1088 -358 1136 -357
rect 1092 -362 1098 -358
rect 1102 -362 1110 -358
rect 1114 -362 1122 -358
rect 1126 -362 1132 -358
rect 780 -389 963 -385
rect 970 -389 1069 -385
rect 137 -689 142 -685
rect 146 -689 154 -685
rect 158 -689 165 -685
rect 169 -689 186 -685
rect 780 -687 784 -389
rect 931 -426 935 -389
rect 970 -394 974 -389
rect 962 -410 966 -404
rect 962 -414 974 -410
rect 1150 -426 1154 -330
rect 1337 -328 1349 -318
rect 1325 -332 1329 -328
rect 1360 -332 1364 -328
rect 1393 -332 1397 -328
rect 1425 -332 1429 -328
rect 1329 -336 1360 -332
rect 1364 -336 1369 -332
rect 1373 -336 1380 -332
rect 1384 -336 1393 -332
rect 1397 -336 1403 -332
rect 1407 -336 1413 -332
rect 1417 -336 1425 -332
rect 1429 -336 1437 -332
rect 931 -430 1154 -426
rect 133 -693 137 -689
rect 72 -727 78 -721
rect 74 -761 78 -727
rect 182 -729 186 -689
rect 540 -691 784 -687
rect 165 -760 169 -753
rect 190 -760 194 -749
rect 540 -760 544 -691
rect 74 -765 133 -761
rect 165 -764 183 -760
rect 190 -764 544 -760
rect 891 -726 1121 -722
rect 80 -772 145 -768
rect 80 -786 84 -772
rect -80 -787 -50 -786
rect -171 -865 -167 -788
rect -68 -790 -50 -787
rect -43 -790 84 -786
rect 98 -779 157 -775
rect -118 -797 -77 -793
rect -118 -799 -114 -797
rect -137 -805 -114 -799
rect -68 -801 -64 -790
rect -43 -795 -39 -790
rect -51 -811 -47 -805
rect -88 -826 -84 -821
rect -51 -826 -38 -811
rect -94 -830 -88 -826
rect -84 -830 -78 -826
rect -74 -830 -68 -826
rect -64 -830 -46 -826
rect -42 -830 -38 -826
rect 13 -837 69 -835
rect 13 -841 15 -837
rect 19 -841 23 -837
rect 27 -841 31 -837
rect 35 -841 50 -837
rect 54 -841 69 -837
rect 13 -843 37 -841
rect 13 -848 17 -843
rect 33 -848 37 -843
rect -288 -870 -6 -865
rect 50 -847 54 -841
rect -339 -878 -295 -874
rect -433 -901 -429 -890
rect -327 -885 -307 -881
rect -474 -905 -440 -901
rect -433 -905 -362 -901
rect -474 -940 -469 -905
rect -433 -910 -429 -905
rect -441 -926 -437 -920
rect -441 -930 -429 -926
rect -327 -940 -322 -885
rect -288 -888 -280 -870
rect -261 -878 -241 -874
rect -11 -876 -6 -870
rect 21 -875 29 -868
rect -11 -880 13 -876
rect 21 -878 37 -875
rect 58 -878 62 -867
rect 98 -876 103 -779
rect 165 -782 169 -764
rect 190 -769 194 -764
rect 141 -786 169 -782
rect 141 -789 149 -786
rect 165 -789 169 -786
rect 891 -778 895 -726
rect 915 -741 941 -736
rect 922 -747 926 -741
rect 930 -778 934 -767
rect 1054 -752 1060 -748
rect 1064 -752 1072 -748
rect 1076 -752 1083 -748
rect 1087 -752 1094 -748
rect 1050 -753 1098 -752
rect 1050 -757 1054 -753
rect 1094 -757 1098 -753
rect 182 -785 186 -779
rect 625 -782 923 -778
rect 930 -782 1038 -778
rect 625 -784 878 -782
rect 182 -789 194 -785
rect 930 -787 934 -782
rect 1012 -785 1019 -782
rect 133 -804 137 -799
rect 153 -804 161 -799
rect 922 -803 926 -797
rect 133 -805 169 -804
rect 137 -809 143 -805
rect 147 -809 155 -805
rect 159 -809 165 -805
rect 922 -807 934 -803
rect 1034 -804 1038 -782
rect 1034 -808 1051 -804
rect 983 -815 1063 -811
rect 983 -831 987 -815
rect 1070 -819 1078 -797
rect 1117 -804 1121 -726
rect 1523 -780 1527 -256
rect 1303 -783 1527 -780
rect 1085 -808 1121 -804
rect 1147 -811 1152 -808
rect 1097 -815 1152 -811
rect 1070 -824 1291 -819
rect 893 -835 987 -831
rect 1019 -832 1063 -828
rect 98 -878 109 -876
rect 21 -879 51 -878
rect -273 -885 -251 -881
rect 33 -882 51 -879
rect 58 -882 109 -878
rect -308 -912 -304 -908
rect -264 -912 -260 -908
rect -308 -913 -260 -912
rect -304 -917 -298 -913
rect -294 -917 -286 -913
rect -282 -917 -274 -913
rect -270 -917 -264 -913
rect -474 -944 -322 -940
rect -254 -951 -251 -885
rect -37 -889 24 -885
rect -351 -960 -238 -951
rect -715 -984 -634 -980
rect -715 -1048 -711 -984
rect -683 -1017 -677 -1013
rect -673 -1017 -667 -1013
rect -663 -1017 -647 -1013
rect -643 -1017 -619 -1013
rect -615 -1017 -587 -1013
rect -583 -1017 -569 -1013
rect -687 -1021 -683 -1017
rect -652 -1021 -648 -1017
rect -619 -1021 -615 -1017
rect -587 -1021 -583 -1017
rect -640 -1041 -628 -1021
rect -607 -1041 -595 -1021
rect -715 -1052 -674 -1048
rect -667 -1049 -663 -1041
rect -632 -1049 -628 -1041
rect -599 -1049 -595 -1041
rect -579 -1049 -575 -1041
rect -715 -1143 -711 -1052
rect -667 -1053 -639 -1049
rect -632 -1053 -618 -1049
rect -599 -1053 -586 -1049
rect -579 -1053 -171 -1049
rect -693 -1059 -686 -1055
rect -667 -1062 -663 -1053
rect -632 -1062 -628 -1053
rect -599 -1062 -595 -1053
rect -579 -1062 -575 -1053
rect -675 -1072 -663 -1062
rect -172 -1055 -171 -1053
rect -172 -1056 -164 -1055
rect -687 -1076 -683 -1072
rect -652 -1076 -648 -1072
rect -619 -1076 -615 -1072
rect -587 -1076 -583 -1072
rect -683 -1080 -652 -1076
rect -648 -1080 -643 -1076
rect -639 -1080 -632 -1076
rect -628 -1080 -619 -1076
rect -615 -1080 -609 -1076
rect -605 -1080 -599 -1076
rect -595 -1080 -587 -1076
rect -583 -1080 -575 -1076
rect -446 -1106 -420 -1101
rect -439 -1112 -435 -1106
rect -431 -1143 -427 -1132
rect -715 -1147 -623 -1143
rect -627 -1191 -623 -1147
rect -473 -1147 -438 -1143
rect -431 -1147 -230 -1143
rect -601 -1160 -595 -1156
rect -591 -1160 -585 -1156
rect -581 -1160 -565 -1156
rect -561 -1160 -537 -1156
rect -533 -1160 -505 -1156
rect -501 -1160 -487 -1156
rect -605 -1164 -601 -1160
rect -570 -1164 -566 -1160
rect -537 -1164 -533 -1160
rect -505 -1164 -501 -1160
rect -558 -1184 -546 -1164
rect -525 -1184 -513 -1164
rect -627 -1195 -592 -1191
rect -585 -1192 -581 -1184
rect -550 -1192 -546 -1184
rect -517 -1192 -513 -1184
rect -497 -1192 -493 -1184
rect -473 -1192 -468 -1147
rect -431 -1152 -427 -1147
rect -439 -1168 -435 -1162
rect -439 -1172 -427 -1168
rect -384 -1170 -328 -1168
rect -627 -1301 -623 -1195
rect -585 -1196 -557 -1192
rect -550 -1196 -536 -1192
rect -517 -1196 -504 -1192
rect -497 -1196 -468 -1192
rect -611 -1202 -604 -1198
rect -585 -1205 -581 -1196
rect -550 -1205 -546 -1196
rect -517 -1205 -513 -1196
rect -497 -1205 -493 -1196
rect -593 -1215 -581 -1205
rect -473 -1206 -468 -1196
rect -384 -1174 -382 -1170
rect -378 -1174 -374 -1170
rect -370 -1174 -366 -1170
rect -362 -1174 -347 -1170
rect -343 -1174 -328 -1170
rect -384 -1176 -360 -1174
rect -384 -1181 -380 -1176
rect -364 -1181 -360 -1176
rect -347 -1180 -343 -1174
rect -473 -1213 -437 -1206
rect -430 -1209 -425 -1206
rect -376 -1208 -368 -1201
rect -430 -1213 -384 -1209
rect -376 -1211 -360 -1208
rect -339 -1211 -335 -1200
rect -376 -1212 -346 -1211
rect -364 -1215 -346 -1212
rect -339 -1215 -322 -1211
rect -605 -1219 -601 -1215
rect -570 -1219 -566 -1215
rect -537 -1219 -533 -1215
rect -505 -1219 -501 -1215
rect -601 -1223 -570 -1219
rect -566 -1223 -561 -1219
rect -557 -1223 -550 -1219
rect -546 -1223 -537 -1219
rect -533 -1223 -527 -1219
rect -523 -1223 -517 -1219
rect -513 -1223 -505 -1219
rect -501 -1223 -493 -1219
rect -472 -1222 -373 -1218
rect -600 -1270 -594 -1266
rect -590 -1270 -584 -1266
rect -580 -1270 -564 -1266
rect -560 -1270 -536 -1266
rect -532 -1270 -504 -1266
rect -500 -1270 -486 -1266
rect -604 -1274 -600 -1270
rect -569 -1274 -565 -1270
rect -536 -1274 -532 -1270
rect -504 -1274 -500 -1270
rect -472 -1274 -468 -1222
rect -364 -1226 -360 -1215
rect -339 -1220 -335 -1215
rect -347 -1236 -343 -1230
rect -384 -1251 -380 -1246
rect -347 -1251 -334 -1236
rect -390 -1255 -384 -1251
rect -380 -1255 -374 -1251
rect -370 -1255 -364 -1251
rect -360 -1255 -342 -1251
rect -338 -1255 -334 -1251
rect -324 -1241 -246 -1236
rect -324 -1274 -320 -1241
rect -557 -1294 -545 -1274
rect -524 -1294 -512 -1274
rect -627 -1305 -591 -1301
rect -584 -1302 -580 -1294
rect -549 -1302 -545 -1294
rect -516 -1302 -512 -1294
rect -496 -1302 -492 -1294
rect -472 -1278 -320 -1274
rect -303 -1252 -297 -1248
rect -293 -1252 -285 -1248
rect -281 -1252 -274 -1248
rect -270 -1252 -263 -1248
rect -307 -1253 -259 -1252
rect -307 -1257 -303 -1253
rect -263 -1257 -259 -1253
rect -472 -1302 -468 -1278
rect -584 -1306 -556 -1302
rect -549 -1306 -535 -1302
rect -516 -1306 -503 -1302
rect -496 -1306 -468 -1302
rect -610 -1312 -603 -1308
rect -584 -1315 -580 -1306
rect -549 -1315 -545 -1306
rect -516 -1315 -512 -1306
rect -496 -1315 -492 -1306
rect -592 -1325 -580 -1315
rect -604 -1329 -600 -1325
rect -569 -1329 -565 -1325
rect -536 -1329 -532 -1325
rect -504 -1329 -500 -1325
rect -600 -1333 -569 -1329
rect -565 -1333 -560 -1329
rect -556 -1333 -549 -1329
rect -545 -1333 -536 -1329
rect -532 -1333 -526 -1329
rect -522 -1333 -516 -1329
rect -512 -1333 -504 -1329
rect -500 -1333 -492 -1329
rect -473 -1355 -468 -1306
rect -430 -1307 -306 -1304
rect -447 -1318 -421 -1313
rect -440 -1324 -436 -1318
rect -338 -1328 -334 -1307
rect -318 -1308 -306 -1307
rect -306 -1315 -294 -1311
rect -287 -1319 -279 -1297
rect -250 -1304 -246 -1241
rect -272 -1308 -246 -1304
rect -234 -1308 -230 -1147
rect -172 -1191 -168 -1056
rect -115 -1152 -59 -1150
rect -115 -1156 -113 -1152
rect -109 -1156 -105 -1152
rect -101 -1156 -97 -1152
rect -93 -1156 -78 -1152
rect -74 -1156 -59 -1152
rect -115 -1158 -91 -1156
rect -115 -1163 -111 -1158
rect -95 -1163 -91 -1158
rect -78 -1162 -74 -1156
rect -107 -1190 -99 -1183
rect -172 -1195 -115 -1191
rect -107 -1193 -91 -1190
rect -70 -1193 -66 -1182
rect -37 -1193 -33 -889
rect 33 -893 37 -882
rect 58 -887 62 -882
rect 893 -894 897 -835
rect 1035 -839 1051 -835
rect 917 -857 943 -852
rect 924 -863 928 -857
rect 932 -894 936 -883
rect 1035 -894 1039 -839
rect 1070 -842 1078 -824
rect 1097 -832 1127 -828
rect 1085 -839 1116 -835
rect 1050 -866 1054 -862
rect 1094 -866 1098 -862
rect 1050 -867 1098 -866
rect 1054 -871 1060 -867
rect 1064 -871 1072 -867
rect 1076 -871 1084 -867
rect 1088 -871 1094 -867
rect 50 -903 54 -897
rect 836 -898 925 -894
rect 932 -898 1031 -894
rect 836 -899 887 -898
rect 13 -918 17 -913
rect 50 -918 63 -903
rect 7 -922 13 -918
rect 17 -922 23 -918
rect 27 -922 33 -918
rect 37 -922 55 -918
rect 59 -922 63 -918
rect 836 -1038 840 -899
rect 893 -935 897 -898
rect 932 -903 936 -898
rect 924 -919 928 -913
rect 924 -923 936 -919
rect 1112 -935 1116 -839
rect 1286 -847 1291 -824
rect 1303 -840 1306 -783
rect 1332 -809 1338 -805
rect 1342 -809 1348 -805
rect 1352 -809 1368 -805
rect 1372 -809 1396 -805
rect 1400 -809 1428 -805
rect 1432 -809 1446 -805
rect 1328 -813 1332 -809
rect 1363 -813 1367 -809
rect 1396 -813 1400 -809
rect 1428 -813 1432 -809
rect 1375 -833 1387 -813
rect 1408 -833 1420 -813
rect 1303 -844 1341 -840
rect 1348 -841 1352 -833
rect 1383 -841 1387 -833
rect 1416 -841 1420 -833
rect 1436 -841 1440 -833
rect 1348 -845 1376 -841
rect 1383 -845 1397 -841
rect 1416 -845 1429 -841
rect 1436 -845 1446 -841
rect 1286 -851 1329 -847
rect 1348 -854 1352 -845
rect 1383 -854 1387 -845
rect 1416 -854 1420 -845
rect 1436 -854 1440 -845
rect 1340 -864 1352 -854
rect 1328 -868 1332 -864
rect 1363 -868 1367 -864
rect 1396 -868 1400 -864
rect 1428 -868 1432 -864
rect 1332 -872 1363 -868
rect 1367 -872 1372 -868
rect 1376 -872 1383 -868
rect 1387 -872 1396 -868
rect 1400 -872 1406 -868
rect 1410 -872 1416 -868
rect 1420 -872 1428 -868
rect 1432 -872 1440 -868
rect 893 -939 1116 -935
rect -107 -1194 -77 -1193
rect -95 -1197 -77 -1194
rect -70 -1197 -33 -1193
rect -260 -1315 -240 -1311
rect -232 -1315 -230 -1308
rect -173 -1204 -104 -1200
rect -173 -1319 -168 -1204
rect -95 -1208 -91 -1197
rect -70 -1202 -66 -1197
rect -78 -1218 -74 -1212
rect -115 -1233 -111 -1228
rect -78 -1233 -65 -1218
rect -121 -1237 -115 -1233
rect -111 -1237 -105 -1233
rect -101 -1237 -95 -1233
rect -91 -1237 -73 -1233
rect -69 -1237 -65 -1233
rect -37 -1290 -33 -1197
rect 487 -1042 840 -1038
rect 5 -1236 11 -1232
rect 15 -1236 21 -1232
rect 25 -1236 35 -1232
rect 1 -1240 5 -1236
rect 31 -1247 35 -1236
rect 31 -1251 38 -1247
rect 42 -1251 57 -1247
rect 31 -1252 57 -1251
rect 38 -1258 42 -1252
rect 21 -1289 25 -1280
rect 46 -1289 50 -1278
rect 487 -1289 491 -1042
rect 867 -1149 1097 -1145
rect 671 -1201 677 -1200
rect 867 -1201 871 -1149
rect 891 -1164 917 -1159
rect 898 -1170 902 -1164
rect 906 -1201 910 -1190
rect 1030 -1175 1036 -1171
rect 1040 -1175 1048 -1171
rect 1052 -1175 1059 -1171
rect 1063 -1175 1070 -1171
rect 1026 -1176 1074 -1175
rect 1026 -1180 1030 -1176
rect 1070 -1180 1074 -1176
rect 671 -1205 899 -1201
rect 906 -1205 1014 -1201
rect 671 -1206 854 -1205
rect 906 -1210 910 -1205
rect 988 -1208 995 -1205
rect 898 -1226 902 -1220
rect 898 -1230 910 -1226
rect 1010 -1227 1014 -1205
rect 1010 -1231 1027 -1227
rect 959 -1238 1039 -1234
rect 959 -1254 963 -1238
rect 1046 -1242 1054 -1220
rect 1093 -1227 1097 -1149
rect 1523 -1195 1527 -783
rect 1298 -1198 1527 -1195
rect 1061 -1231 1097 -1227
rect 1123 -1234 1128 -1231
rect 1073 -1238 1128 -1234
rect 1046 -1247 1287 -1242
rect -37 -1294 13 -1290
rect 21 -1293 39 -1289
rect 46 -1293 491 -1289
rect 869 -1258 963 -1254
rect 995 -1255 1039 -1251
rect -128 -1297 -127 -1295
rect 21 -1297 25 -1293
rect -128 -1301 1 -1297
rect 9 -1300 25 -1297
rect 46 -1298 50 -1293
rect 9 -1304 17 -1300
rect -287 -1324 -168 -1319
rect 1 -1319 5 -1314
rect 21 -1319 25 -1314
rect 38 -1314 42 -1308
rect 38 -1318 43 -1314
rect 47 -1318 50 -1314
rect 869 -1316 873 -1258
rect 1011 -1262 1027 -1258
rect 893 -1280 919 -1275
rect 900 -1286 904 -1280
rect 758 -1317 873 -1316
rect 908 -1317 912 -1306
rect 1011 -1317 1015 -1262
rect 1046 -1265 1054 -1247
rect 1073 -1255 1103 -1251
rect 1282 -1257 1287 -1247
rect 1298 -1250 1301 -1198
rect 1324 -1219 1330 -1215
rect 1334 -1219 1340 -1215
rect 1344 -1219 1360 -1215
rect 1364 -1219 1388 -1215
rect 1392 -1219 1420 -1215
rect 1424 -1219 1438 -1215
rect 1320 -1223 1324 -1219
rect 1355 -1223 1359 -1219
rect 1388 -1223 1392 -1219
rect 1420 -1223 1424 -1219
rect 1367 -1243 1379 -1223
rect 1400 -1243 1412 -1223
rect 1298 -1254 1333 -1250
rect 1340 -1251 1344 -1243
rect 1375 -1251 1379 -1243
rect 1408 -1251 1412 -1243
rect 1428 -1251 1432 -1243
rect 1340 -1255 1368 -1251
rect 1375 -1255 1389 -1251
rect 1408 -1255 1421 -1251
rect 1428 -1255 1438 -1251
rect 1061 -1262 1092 -1258
rect 1282 -1261 1321 -1257
rect 1026 -1289 1030 -1285
rect 1070 -1289 1074 -1285
rect 1026 -1290 1074 -1289
rect 1030 -1294 1036 -1290
rect 1040 -1294 1048 -1290
rect 1052 -1294 1060 -1290
rect 1064 -1294 1070 -1290
rect 38 -1319 41 -1318
rect 1 -1320 41 -1319
rect 5 -1324 11 -1320
rect 15 -1324 21 -1320
rect 25 -1324 41 -1320
rect 758 -1321 901 -1317
rect 908 -1321 1007 -1317
rect -338 -1332 -294 -1328
rect -432 -1355 -428 -1344
rect -326 -1339 -306 -1335
rect -473 -1359 -439 -1355
rect -432 -1359 -361 -1355
rect -473 -1394 -468 -1359
rect -432 -1364 -428 -1359
rect -440 -1380 -436 -1374
rect -440 -1384 -428 -1380
rect -326 -1394 -321 -1339
rect -287 -1342 -279 -1324
rect -260 -1332 -240 -1328
rect -272 -1339 -250 -1335
rect -307 -1366 -303 -1362
rect -263 -1366 -259 -1362
rect -307 -1367 -259 -1366
rect -303 -1371 -297 -1367
rect -293 -1371 -285 -1367
rect -281 -1371 -273 -1367
rect -269 -1371 -263 -1367
rect -473 -1398 -321 -1394
rect -253 -1405 -250 -1339
rect -193 -1377 -189 -1324
rect 758 -1376 763 -1321
rect 869 -1358 873 -1321
rect 908 -1326 912 -1321
rect 900 -1342 904 -1336
rect 900 -1346 912 -1342
rect 1088 -1358 1092 -1262
rect 1340 -1264 1344 -1255
rect 1375 -1264 1379 -1255
rect 1408 -1264 1412 -1255
rect 1428 -1264 1432 -1255
rect 1332 -1274 1344 -1264
rect 1320 -1278 1324 -1274
rect 1355 -1278 1359 -1274
rect 1388 -1278 1392 -1274
rect 1420 -1278 1424 -1274
rect 1324 -1282 1355 -1278
rect 1359 -1282 1364 -1278
rect 1368 -1282 1375 -1278
rect 1379 -1282 1388 -1278
rect 1392 -1282 1398 -1278
rect 1402 -1282 1408 -1278
rect 1412 -1282 1420 -1278
rect 1424 -1282 1432 -1278
rect 869 -1362 1092 -1358
rect 106 -1377 763 -1376
rect -193 -1381 763 -1377
rect -350 -1414 -237 -1405
<< m2contact >>
rect 1224 923 1231 930
rect 487 883 492 891
rect 338 631 345 637
rect -439 549 -432 556
rect -326 547 -321 553
rect -439 455 -432 462
rect -315 443 -308 451
rect -242 447 -234 454
rect -173 564 -164 569
rect -363 403 -352 410
rect -242 428 -234 434
rect 847 695 852 700
rect 1059 575 1066 582
rect 1168 563 1174 570
rect 1199 552 1206 559
rect -143 377 -138 383
rect -362 348 -352 357
rect 12 378 17 383
rect -439 149 -432 156
rect -326 147 -321 153
rect -439 55 -432 62
rect -315 43 -308 51
rect -242 47 -234 54
rect 115 357 120 362
rect 1059 534 1066 541
rect 58 164 65 170
rect -185 155 -179 161
rect 241 299 246 304
rect 1174 534 1180 540
rect 761 455 768 462
rect 1078 466 1086 473
rect 117 163 128 168
rect 161 164 169 169
rect -363 3 -352 10
rect -242 28 -234 34
rect 163 83 169 88
rect -102 7 -95 14
rect -362 -52 -352 -43
rect -440 -298 -433 -291
rect -312 -300 -306 -294
rect -440 -392 -433 -385
rect -316 -404 -309 -396
rect -243 -400 -235 -393
rect 98 7 105 14
rect 313 223 318 228
rect 228 164 237 169
rect 231 83 238 88
rect 888 184 894 190
rect 1059 175 1066 182
rect 1168 163 1174 170
rect 1199 152 1206 159
rect 468 126 475 133
rect 1059 134 1066 141
rect 1174 134 1180 140
rect 180 -98 186 -92
rect 255 -218 261 -212
rect 228 -253 235 -246
rect -157 -290 -151 -284
rect 1078 66 1086 73
rect -57 -362 -51 -355
rect -364 -444 -353 -437
rect -243 -419 -235 -413
rect -363 -499 -353 -490
rect -438 -759 -431 -752
rect -317 -761 -311 -755
rect -438 -853 -431 -846
rect -314 -865 -307 -857
rect -241 -861 -233 -854
rect 61 -434 67 -428
rect 228 -432 235 -425
rect 109 -446 115 -439
rect 1050 -283 1057 -276
rect 1159 -295 1165 -288
rect 1190 -306 1197 -299
rect 1050 -324 1057 -317
rect 1165 -324 1171 -318
rect 1069 -392 1077 -385
rect 72 -721 78 -715
rect -143 -805 -137 -799
rect -362 -905 -351 -898
rect -241 -880 -233 -874
rect -48 -876 -42 -870
rect 619 -784 625 -778
rect 1012 -792 1019 -785
rect 1121 -804 1127 -797
rect 1152 -815 1159 -808
rect 1012 -833 1019 -826
rect 109 -882 115 -876
rect -361 -960 -351 -951
rect -171 -1055 -164 -1049
rect -437 -1213 -430 -1206
rect -322 -1215 -316 -1209
rect -437 -1307 -430 -1300
rect -313 -1319 -306 -1311
rect 1127 -833 1133 -827
rect 1031 -901 1039 -894
rect -240 -1315 -232 -1308
rect 665 -1206 671 -1200
rect 988 -1215 995 -1208
rect 1097 -1227 1103 -1220
rect 1128 -1238 1135 -1231
rect 988 -1256 995 -1249
rect -134 -1301 -128 -1295
rect 1103 -1256 1109 -1250
rect -361 -1359 -350 -1352
rect -240 -1334 -232 -1328
rect 1007 -1324 1015 -1317
rect -360 -1414 -350 -1405
<< metal2 >>
rect 1224 890 1231 923
rect 492 883 1231 890
rect -166 766 852 771
rect -166 637 -161 766
rect 847 700 852 766
rect -326 632 338 637
rect -439 462 -432 549
rect -326 553 -321 632
rect -363 440 -308 443
rect -363 410 -352 440
rect -242 434 -234 447
rect -362 357 -352 403
rect -352 348 -351 354
rect -171 237 -166 564
rect 1059 541 1066 575
rect 1174 540 1180 570
rect 1199 473 1206 552
rect 1086 466 1206 473
rect 468 455 761 462
rect -138 378 12 383
rect -63 336 -58 378
rect 75 357 115 362
rect -63 331 -5 336
rect -10 325 -5 331
rect 75 325 80 357
rect -10 320 80 325
rect 59 309 64 320
rect 59 304 205 309
rect 200 299 241 304
rect -326 232 318 237
rect -439 62 -432 149
rect -326 153 -321 232
rect 313 228 318 232
rect 65 164 117 168
rect 128 164 131 168
rect 169 164 228 168
rect -363 40 -308 43
rect -363 10 -352 40
rect -242 34 -234 47
rect -362 -43 -352 3
rect -352 -52 -351 -46
rect -185 -212 -179 155
rect 468 133 475 455
rect 649 184 888 190
rect 169 83 231 87
rect -95 7 98 14
rect 27 -100 33 7
rect 180 -100 186 -98
rect 27 -106 186 -100
rect 27 -162 33 -106
rect 649 -162 655 184
rect 1059 141 1066 175
rect 1174 140 1180 170
rect 1199 73 1206 152
rect 1086 66 1206 73
rect 27 -168 655 -162
rect -312 -218 255 -212
rect -440 -385 -433 -298
rect -312 -294 -306 -218
rect -364 -407 -309 -404
rect -364 -437 -353 -407
rect -243 -413 -235 -400
rect -363 -490 -353 -444
rect -353 -499 -352 -493
rect -157 -715 -151 -290
rect -57 -428 -51 -362
rect 228 -425 235 -253
rect 1050 -317 1057 -283
rect 1165 -318 1171 -288
rect 1190 -385 1197 -306
rect 1077 -392 1197 -385
rect -57 -434 61 -428
rect -317 -721 72 -715
rect -438 -846 -431 -759
rect -317 -755 -311 -721
rect -362 -868 -307 -865
rect -362 -898 -351 -868
rect -241 -874 -233 -861
rect -361 -951 -351 -905
rect -351 -960 -350 -954
rect -143 -1025 -137 -805
rect -48 -936 -42 -876
rect 109 -876 115 -446
rect 619 -936 625 -784
rect 1012 -826 1019 -792
rect 1127 -827 1133 -797
rect 1152 -894 1159 -815
rect 1039 -901 1159 -894
rect -48 -942 625 -936
rect -220 -1031 -137 -1025
rect -220 -1209 -214 -1031
rect -164 -1055 -131 -1049
rect -137 -1125 -131 -1055
rect -137 -1131 671 -1125
rect 665 -1200 671 -1131
rect -437 -1300 -430 -1213
rect -316 -1215 -214 -1209
rect -220 -1280 -214 -1215
rect 988 -1249 995 -1215
rect 1103 -1250 1109 -1220
rect -220 -1286 -128 -1280
rect -134 -1295 -128 -1286
rect -134 -1302 -128 -1301
rect -361 -1322 -306 -1319
rect -361 -1352 -350 -1322
rect -240 -1328 -232 -1315
rect 1128 -1317 1135 -1238
rect 1015 -1324 1135 -1317
rect -360 -1405 -350 -1359
rect -350 -1414 -349 -1408
<< labels >>
rlabel metal1 915 -741 941 -736 5 vdd
rlabel metal1 925 -806 930 -805 1 gnd
rlabel metal1 917 -857 943 -852 5 vdd
rlabel metal1 927 -922 932 -921 1 gnd
rlabel metal1 1078 -751 1081 -749 5 vdd
rlabel metal1 1078 -870 1081 -868 1 gnd
rlabel metal1 953 -232 979 -227 5 vdd
rlabel metal1 963 -297 968 -296 1 gnd
rlabel metal1 955 -348 981 -343 5 vdd
rlabel metal1 965 -413 970 -412 1 gnd
rlabel metal1 1116 -242 1119 -240 5 vdd
rlabel metal1 1116 -361 1119 -359 1 gnd
rlabel metal1 962 226 988 231 5 vdd
rlabel metal1 972 161 977 162 1 gnd
rlabel metal1 964 110 990 115 5 vdd
rlabel metal1 974 45 979 46 1 gnd
rlabel metal1 1125 216 1128 218 5 vdd
rlabel metal1 1125 97 1128 99 1 gnd
rlabel metal1 1213 144 1216 147 7 s3
rlabel metal1 1204 -314 1207 -311 1 s2
rlabel metal1 1166 -823 1169 -820 1 s1
rlabel metal1 1323 -843 1325 -841 3 clk
rlabel metal1 1390 -871 1392 -869 1 gnd
rlabel metal1 1390 -808 1392 -806 5 vdd
rlabel metal1 1375 -808 1377 -806 5 vdd
rlabel metal1 1334 -808 1336 -806 5 vdd
rlabel metal1 1335 -871 1337 -869 1 gnd
rlabel metal1 1434 -871 1436 -869 1 gnd
rlabel metal1 1434 -808 1436 -806 5 vdd
rlabel metal1 1441 -844 1444 -842 1 s1q
rlabel metal1 1320 -307 1322 -305 3 clk
rlabel metal1 1387 -335 1389 -333 1 gnd
rlabel metal1 1387 -272 1389 -270 5 vdd
rlabel metal1 1372 -272 1374 -270 5 vdd
rlabel metal1 1331 -272 1333 -270 5 vdd
rlabel metal1 1332 -335 1334 -333 1 gnd
rlabel metal1 1431 -335 1433 -333 1 gnd
rlabel metal1 1431 -272 1433 -270 5 vdd
rlabel metal1 1439 -308 1441 -305 1 s2q
rlabel metal1 1323 154 1325 156 3 clk
rlabel metal1 1390 126 1392 128 1 gnd
rlabel metal1 1390 189 1392 191 5 vdd
rlabel metal1 1375 189 1377 191 5 vdd
rlabel metal1 1334 189 1336 191 5 vdd
rlabel metal1 1335 126 1337 128 1 gnd
rlabel metal1 1434 126 1436 128 1 gnd
rlabel metal1 1434 189 1436 191 5 vdd
rlabel metal1 1442 153 1444 155 1 s3q
rlabel metal1 1434 -1254 1437 -1252 1 s0q
rlabel metal1 1426 -1218 1428 -1216 5 vdd
rlabel metal1 1426 -1281 1428 -1279 1 gnd
rlabel metal1 1327 -1281 1329 -1279 1 gnd
rlabel metal1 1326 -1218 1328 -1216 5 vdd
rlabel metal1 1367 -1218 1369 -1216 5 vdd
rlabel metal1 1382 -1218 1384 -1216 5 vdd
rlabel metal1 1382 -1281 1384 -1279 1 gnd
rlabel metal1 1315 -1253 1317 -1251 3 clk
rlabel metal1 1143 -1246 1146 -1243 1 s0
rlabel metal1 1054 -1293 1057 -1291 1 gnd
rlabel metal1 1054 -1174 1057 -1172 5 vdd
rlabel metal1 903 -1345 908 -1344 1 gnd
rlabel metal1 893 -1280 919 -1275 5 vdd
rlabel metal1 901 -1229 906 -1228 1 gnd
rlabel metal1 891 -1164 917 -1159 5 vdd
rlabel metal1 450 127 452 129 7 c4
rlabel metal1 391 267 394 269 5 vdd
rlabel metal1 391 91 394 93 1 gnd
rlabel metal1 307 -99 309 -97 1 p3p2p1p0c0
rlabel metal1 296 -124 301 -123 1 gnd
rlabel metal1 286 -59 312 -54 5 vdd
rlabel metal1 267 -61 269 -60 1 vdd
rlabel metal1 180 -12 182 -10 1 p3p2p1g0
rlabel metal1 168 -37 173 -36 1 gnd
rlabel metal1 158 28 184 33 5 vdd
rlabel metal1 139 26 141 27 1 vdd
rlabel metal1 64 84 66 86 1 p3p2g1
rlabel metal1 53 59 58 60 1 gnd
rlabel metal1 43 124 69 129 5 vdd
rlabel metal1 24 122 26 123 1 vdd
rlabel metal1 -55 165 -53 167 1 p3g2
rlabel metal1 -66 140 -61 141 1 gnd
rlabel metal1 -76 205 -50 210 5 vdd
rlabel metal1 -95 203 -93 204 1 vdd
rlabel metal1 385 -296 387 -294 7 c3
rlabel metal1 337 -339 339 -337 1 gnd
rlabel metal1 336 -198 338 -196 5 vdd
rlabel metal1 217 -435 219 -433 7 p2p1p0c0
rlabel metal1 205 -460 210 -459 1 gnd
rlabel metal1 195 -395 221 -390 5 vdd
rlabel metal1 176 -397 178 -396 1 vdd
rlabel metal1 65 -881 68 -879 1 p1p0c0
rlabel metal1 73 -353 75 -350 1 p2p1g0
rlabel metal1 62 -377 67 -376 1 gnd
rlabel metal1 52 -312 78 -307 5 vdd
rlabel metal1 33 -314 35 -313 1 vdd
rlabel metal1 -57 -280 -55 -278 1 p2g1
rlabel metal1 -69 -305 -64 -304 1 gnd
rlabel metal1 -79 -240 -53 -235 5 vdd
rlabel metal1 -98 -242 -96 -241 1 vdd
rlabel metal1 196 -763 199 -761 7 c2
rlabel metal1 149 -808 151 -806 1 gnd
rlabel metal1 148 -688 151 -686 5 vdd
rlabel metal1 185 -788 190 -787 1 gnd
rlabel metal1 -36 -789 -34 -787 1 p1g0
rlabel metal1 -48 -814 -43 -813 1 gnd
rlabel metal1 -58 -749 -32 -744 5 vdd
rlabel metal1 -77 -751 -75 -750 1 vdd
rlabel metal1 53 -906 58 -905 1 gnd
rlabel metal1 43 -841 69 -836 5 vdd
rlabel metal1 24 -843 26 -842 1 vdd
rlabel metal1 53 -1292 55 -1290 7 c1
rlabel metal1 17 -1235 19 -1233 1 vdd
rlabel metal1 17 -1323 19 -1321 1 gnd
rlabel metal1 -63 -1196 -60 -1194 7 p0c0
rlabel metal1 -75 -1221 -70 -1220 1 gnd
rlabel metal1 -85 -1156 -59 -1151 5 vdd
rlabel metal1 -104 -1158 -102 -1157 1 vdd
rlabel metal1 -573 -1052 -571 -1050 7 c0
rlabel metal1 -692 -1058 -690 -1056 1 c0d
rlabel metal1 -581 -1016 -579 -1014 5 vdd
rlabel metal1 -581 -1079 -579 -1077 1 gnd
rlabel metal1 -680 -1079 -678 -1077 1 gnd
rlabel metal1 -681 -1016 -679 -1014 5 vdd
rlabel metal1 -640 -1016 -638 -1014 5 vdd
rlabel metal1 -625 -1016 -623 -1014 5 vdd
rlabel metal1 -625 -1079 -623 -1077 1 gnd
rlabel metal1 -692 -1051 -690 -1049 3 clk
rlabel metal1 -492 -386 -490 -384 1 b2
rlabel metal1 -611 -392 -609 -390 1 b2d
rlabel metal1 -500 -350 -498 -348 5 vdd
rlabel metal1 -500 -413 -498 -411 1 gnd
rlabel metal1 -599 -413 -597 -411 1 gnd
rlabel metal1 -600 -350 -598 -348 5 vdd
rlabel metal1 -559 -350 -557 -348 5 vdd
rlabel metal1 -544 -350 -542 -348 5 vdd
rlabel metal1 -544 -413 -542 -411 1 gnd
rlabel metal1 -611 -385 -609 -383 3 clk
rlabel metal1 -612 -751 -610 -749 1 a1d
rlabel metal1 -493 -745 -491 -743 1 a1
rlabel metal1 -501 -709 -499 -707 5 vdd
rlabel metal1 -501 -772 -499 -770 1 gnd
rlabel metal1 -600 -772 -598 -770 1 gnd
rlabel metal1 -601 -709 -599 -707 5 vdd
rlabel metal1 -560 -709 -558 -707 5 vdd
rlabel metal1 -545 -709 -543 -707 5 vdd
rlabel metal1 -545 -772 -543 -770 1 gnd
rlabel metal1 -612 -744 -610 -742 3 clk
rlabel metal1 -491 -848 -489 -846 7 b1
rlabel metal1 -610 -854 -608 -852 1 b1d
rlabel metal1 -499 -812 -497 -810 5 vdd
rlabel metal1 -499 -875 -497 -873 1 gnd
rlabel metal1 -598 -875 -596 -873 1 gnd
rlabel metal1 -599 -812 -597 -810 5 vdd
rlabel metal1 -558 -812 -556 -810 5 vdd
rlabel metal1 -543 -812 -541 -810 5 vdd
rlabel metal1 -543 -875 -541 -873 1 gnd
rlabel metal1 -610 -847 -608 -845 3 clk
rlabel metal1 -610 -1201 -608 -1199 3 a0d
rlabel metal1 -423 -1359 -419 -1355 1 b0bar
rlabel metal1 -422 -1147 -418 -1143 1 a0bar
rlabel metal1 -332 -1215 -328 -1211 1 g0
rlabel metal1 -217 -1323 -214 -1320 7 p0
rlabel metal1 -279 -1370 -276 -1368 1 gnd
rlabel metal1 -279 -1251 -276 -1249 5 vdd
rlabel metal1 -344 -1239 -339 -1238 1 gnd
rlabel metal1 -354 -1174 -328 -1169 5 vdd
rlabel metal1 -373 -1176 -371 -1175 1 vdd
rlabel metal1 -437 -1383 -432 -1382 1 gnd
rlabel metal1 -447 -1318 -421 -1313 5 vdd
rlabel metal1 -436 -1171 -431 -1170 1 gnd
rlabel metal1 -446 -1106 -420 -1101 5 vdd
rlabel metal1 -424 -904 -421 -901 1 b1bar
rlabel metal1 -423 -693 -420 -690 1 a1bar
rlabel metal1 -333 -761 -329 -757 1 g1
rlabel metal1 -218 -869 -216 -867 7 p1
rlabel metal1 -280 -916 -277 -914 1 gnd
rlabel metal1 -280 -797 -277 -795 5 vdd
rlabel metal1 -345 -785 -340 -784 1 gnd
rlabel metal1 -355 -720 -329 -715 5 vdd
rlabel metal1 -374 -722 -372 -721 1 vdd
rlabel metal1 -438 -929 -433 -928 1 gnd
rlabel metal1 -448 -864 -422 -859 5 vdd
rlabel metal1 -437 -717 -432 -716 1 gnd
rlabel metal1 -447 -652 -421 -647 5 vdd
rlabel metal1 -609 -1311 -607 -1309 1 b0d
rlabel metal1 -490 -1305 -488 -1303 7 b0
rlabel metal1 -491 -1195 -489 -1193 7 a0
rlabel metal1 -498 -1269 -496 -1267 5 vdd
rlabel metal1 -498 -1332 -496 -1330 1 gnd
rlabel metal1 -597 -1332 -595 -1330 1 gnd
rlabel metal1 -598 -1269 -596 -1267 5 vdd
rlabel metal1 -557 -1269 -555 -1267 5 vdd
rlabel metal1 -542 -1269 -540 -1267 5 vdd
rlabel metal1 -542 -1332 -540 -1330 1 gnd
rlabel metal1 -609 -1304 -607 -1302 3 clk
rlabel metal1 -499 -1159 -497 -1157 5 vdd
rlabel metal1 -499 -1222 -497 -1220 1 gnd
rlabel metal1 -598 -1222 -596 -1220 1 gnd
rlabel metal1 -599 -1159 -597 -1157 5 vdd
rlabel metal1 -558 -1159 -556 -1157 5 vdd
rlabel metal1 -543 -1159 -541 -1157 5 vdd
rlabel metal1 -543 -1222 -541 -1220 1 gnd
rlabel metal1 -610 -1194 -608 -1192 3 clk
rlabel metal1 -426 -443 -423 -440 1 b2bar
rlabel metal1 -425 -232 -422 -229 1 a2bar
rlabel metal1 -335 -299 -332 -296 1 g2
rlabel metal1 -218 -408 -215 -405 7 p2
rlabel metal1 -282 -455 -279 -453 1 gnd
rlabel metal1 -282 -336 -279 -334 5 vdd
rlabel metal1 -347 -324 -342 -323 1 gnd
rlabel metal1 -357 -259 -331 -254 5 vdd
rlabel metal1 -376 -261 -374 -260 1 vdd
rlabel metal1 -440 -468 -435 -467 1 gnd
rlabel metal1 -450 -403 -424 -398 5 vdd
rlabel metal1 -439 -256 -434 -255 1 gnd
rlabel metal1 -449 -191 -423 -186 5 vdd
rlabel metal1 -491 -284 -489 -282 7 a2
rlabel metal1 -610 -290 -608 -288 1 a2d
rlabel metal1 -499 -248 -497 -246 5 vdd
rlabel metal1 -499 -311 -497 -309 1 gnd
rlabel metal1 -598 -311 -596 -309 1 gnd
rlabel metal1 -599 -248 -597 -246 5 vdd
rlabel metal1 -558 -248 -556 -246 5 vdd
rlabel metal1 -543 -248 -541 -246 5 vdd
rlabel metal1 -543 -311 -541 -309 1 gnd
rlabel metal1 -610 -283 -608 -281 3 clk
rlabel metal1 -217 39 -214 42 7 p3
rlabel metal1 -281 -8 -278 -6 1 gnd
rlabel metal1 -281 111 -278 113 5 vdd
rlabel metal1 -334 148 -332 150 7 g3
rlabel metal1 -346 123 -341 124 1 gnd
rlabel metal1 -356 188 -330 193 5 vdd
rlabel metal1 -375 186 -373 187 1 vdd
rlabel metal1 -425 4 -423 6 7 b3bar
rlabel metal1 -423 216 -421 218 7 a3bar
rlabel metal1 -439 -21 -434 -20 1 gnd
rlabel metal1 -449 44 -423 49 5 vdd
rlabel metal1 -438 191 -433 192 1 gnd
rlabel metal1 -448 256 -422 261 5 vdd
rlabel metal1 -491 61 -489 63 7 b3
rlabel metal1 -608 157 -606 159 1 a3d
rlabel metal1 -610 55 -608 57 1 b3d
rlabel metal1 -499 97 -497 99 5 vdd
rlabel metal1 -499 34 -497 36 1 gnd
rlabel metal1 -598 34 -596 36 1 gnd
rlabel metal1 -599 97 -597 99 5 vdd
rlabel metal1 -558 97 -556 99 5 vdd
rlabel metal1 -543 97 -541 99 5 vdd
rlabel metal1 -543 34 -541 36 1 gnd
rlabel metal1 -610 62 -608 64 3 clk
rlabel metal1 -489 163 -487 165 7 a3
rlabel metal1 -497 199 -495 201 5 vdd
rlabel metal1 -497 136 -495 138 1 gnd
rlabel metal1 -596 136 -594 138 1 gnd
rlabel metal1 -597 199 -595 201 5 vdd
rlabel metal1 -556 199 -554 201 5 vdd
rlabel metal1 -541 199 -539 201 5 vdd
rlabel metal1 -541 136 -539 138 1 gnd
rlabel metal1 -608 164 -606 166 3 clk
rlabel metal1 1329 940 1331 942 3 clk
rlabel metal1 1396 912 1398 914 1 gnd
rlabel metal1 1396 975 1398 977 5 vdd
rlabel metal1 1381 975 1383 977 5 vdd
rlabel metal1 1340 975 1342 977 5 vdd
rlabel metal1 1341 912 1343 914 1 gnd
rlabel metal1 1440 912 1442 914 1 gnd
rlabel metal1 1440 975 1442 977 5 vdd
rlabel metal1 -608 564 -606 566 3 clk
rlabel metal1 -541 536 -539 538 1 gnd
rlabel metal1 -541 599 -539 601 5 vdd
rlabel metal1 -556 599 -554 601 5 vdd
rlabel metal1 -597 599 -595 601 5 vdd
rlabel metal1 -596 536 -594 538 1 gnd
rlabel metal1 -497 536 -495 538 1 gnd
rlabel metal1 -497 599 -495 601 5 vdd
rlabel metal1 -610 462 -608 464 3 clk
rlabel metal1 -543 434 -541 436 1 gnd
rlabel metal1 -543 497 -541 499 5 vdd
rlabel metal1 -558 497 -556 499 5 vdd
rlabel metal1 -599 497 -597 499 5 vdd
rlabel metal1 -598 434 -596 436 1 gnd
rlabel metal1 -499 434 -497 436 1 gnd
rlabel metal1 -499 497 -497 499 5 vdd
rlabel metal1 -448 656 -422 661 5 vdd
rlabel metal1 -438 591 -433 592 1 gnd
rlabel metal1 -449 444 -423 449 5 vdd
rlabel metal1 -439 379 -434 380 1 gnd
rlabel metal1 -375 586 -373 587 1 vdd
rlabel metal1 -356 588 -330 593 5 vdd
rlabel metal1 -346 523 -341 524 1 gnd
rlabel metal1 -281 511 -278 513 5 vdd
rlabel metal1 -281 392 -278 394 1 gnd
rlabel metal1 962 626 988 631 5 vdd
rlabel metal1 972 561 977 562 1 gnd
rlabel metal1 964 510 990 515 5 vdd
rlabel metal1 974 445 979 446 1 gnd
rlabel metal1 1125 616 1128 618 5 vdd
rlabel metal1 1125 497 1128 499 1 gnd
rlabel metal1 1323 554 1325 556 3 clk
rlabel metal1 1390 526 1392 528 1 gnd
rlabel metal1 1390 589 1392 591 5 vdd
rlabel metal1 1375 589 1377 591 5 vdd
rlabel metal1 1334 589 1336 591 5 vdd
rlabel metal1 1335 526 1337 528 1 gnd
rlabel metal1 1434 526 1436 528 1 gnd
rlabel metal1 1434 589 1436 591 5 vdd
rlabel metal1 -610 455 -608 457 1 b4d
rlabel metal1 -608 557 -606 559 1 a4d
rlabel metal1 -491 461 -489 463 1 b4
rlabel metal1 -489 563 -487 565 1 a4
rlabel metal1 -423 616 -421 618 1 a4-bar
rlabel metal1 -425 404 -423 406 1 b4-bar
rlabel metal1 -334 548 -332 550 1 g4
rlabel metal1 -217 439 -214 442 1 p4
rlabel metal1 448 529 450 531 1 nout
rlabel metal1 387 551 390 553 3 e
rlabel metal1 387 544 390 546 3 d
rlabel metal1 387 537 390 539 3 c
rlabel metal1 387 530 390 532 3 b
rlabel metal1 387 523 390 525 3 a
rlabel metal1 419 493 422 495 1 gnd
rlabel metal1 369 560 371 562 3 f
rlabel metal1 478 540 483 541 1 c5
rlabel metal1 -128 610 -126 611 1 vdd
rlabel metal1 -143 574 -141 576 3 b
rlabel metal1 -143 565 -141 567 3 a
rlabel metal1 -118 567 -116 569 1 nout
rlabel metal1 -109 612 -83 617 5 vdd
rlabel metal1 -99 547 -94 548 1 gnd
rlabel metal1 1213 544 1216 547 1 s4
rlabel metal1 1442 553 1444 555 1 s4d
rlabel metal1 -88 573 -83 574 1 p4g3
rlabel metal1 -55 516 -53 517 1 vdd
rlabel metal1 -70 480 -68 482 3 b
rlabel metal1 -70 471 -68 473 3 a
rlabel metal1 -45 473 -43 475 1 nout
rlabel metal1 -36 518 -10 523 5 vdd
rlabel metal1 -15 479 -10 480 7 out
rlabel metal1 -26 453 -21 454 1 gnd
rlabel metal1 -17 478 -13 480 1 p4p3g2
rlabel metal1 31 415 33 416 1 vdd
rlabel metal1 16 379 18 381 3 b
rlabel metal1 16 370 18 372 3 a
rlabel metal1 41 372 43 374 1 nout
rlabel metal1 50 417 76 422 5 vdd
rlabel metal1 60 352 65 353 1 gnd
rlabel metal1 69 376 76 380 1 p4p3p2g1
rlabel metal1 136 395 138 396 1 vdd
rlabel metal1 121 359 123 361 3 b
rlabel metal1 121 350 123 352 3 a
rlabel metal1 146 352 148 354 1 nout
rlabel metal1 155 397 181 402 5 vdd
rlabel metal1 165 332 170 333 1 gnd
rlabel metal1 174 357 181 359 1 p4p3p2p1g0
rlabel metal1 262 336 264 337 1 vdd
rlabel metal1 247 300 249 302 3 b
rlabel metal1 247 291 249 293 3 a
rlabel metal1 272 293 274 295 1 nout
rlabel metal1 281 338 307 343 5 vdd
rlabel metal1 291 273 296 274 1 gnd
rlabel metal1 300 297 307 301 1 p4p3p2p1p0g0
rlabel metal1 1448 939 1451 942 1 c5d
rlabel metal1 419 706 422 708 5 vdd
<< end >>
