.include TSMC_180nm.txt
.param SUPPLY=1.8
.option scale=90n
.global gnd vdd

Vdd vdd gnd 'SUPPLY'

M1000 a_n6_n23# a vdd vdd CMOSP w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=90u
M1001 nout b a_n6_n23# vdd CMOSP w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=50u
M1002 out nout vdd vdd CMOSP w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1003 gnd b nout Gnd CMOSN w=10 l=2
+  ad=50p pd=30u as=50p ps=20u
M1004 nout a gnd Gnd CMOSN w=10 l=2
+  ad=50p pd=20u as=50p ps=30u
M1005 out nout gnd Gnd CMOSN w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
C0 nout gnd 0.34799f
C1 a gnd 0.056598f
C2 vdd nout 0.113211f
C3 vdd a 0.020635f
C4 out gnd 0.123714f
C5 b gnd 0.001614f
C6 vdd out 0.243018f
C7 a nout 0.057525f
C8 vdd b 0.020182f
C9 nout out 0.060313f
C10 b nout 0.190775f
C11 vdd a_n6_n23# 1.36e-19
C12 a b 0.190682f
C13 gnd 0 0.237274f 
C14 out 0 0.106495f 
C15 nout 0 0.398928f 
C16 b 0 0.266055f 
C17 a 0 0.230766f 
C18 vdd 0 3.9854f 


va a gnd pulse 0 1.8 0 0.1n 0.1n 10n 20n
vb b gnd pulse 0 1.8 0 0.1n 0.1n 20n 40n

* Propagation delay measurements: input (a,b) -> out
.measure tran tpd_a_lh TRIG v(a) VAL=0.9 RISE=1 TARG v(out) VAL=0.9 RISE=1
.measure tran tpd_a_hl TRIG v(a) VAL=0.9 RISE=2 TARG v(out) VAL=0.9 FALL=1
.measure tran avg_tpd_a param = ((tpd_a_lh + tpd_a_hl)/2)

.measure tran tpd_b_lh TRIG v(b) VAL=0.9 RISE=1 TARG v(out) VAL=0.9 RISE=1
.measure tran tpd_b_hl TRIG v(b) VAL=0.9 RISE=2 TARG v(out) VAL=0.9 FALL=1
.measure tran avg_tpd_b param = ((tpd_b_lh + tpd_b_hl)/2)

.tran  0.01n 100ns
.control
run
plot v(a) v(b)+2 v(out)+4
set hcopypscolor = 1
set color0=white
set color1=black
.endc