magic
tech scmos
timestamp 1731330865
<< nwell >>
rect -9 -5 17 29
<< ntransistor >>
rect 3 -28 5 -18
<< ptransistor >>
rect 3 2 5 22
<< ndiffusion >>
rect 2 -28 3 -18
rect 5 -28 6 -18
<< pdiffusion >>
rect 2 2 3 22
rect 5 2 6 22
<< ndcontact >>
rect -2 -28 2 -18
rect 6 -28 10 -18
<< pdcontact >>
rect -2 2 2 22
rect 6 2 10 22
<< polysilicon >>
rect 3 22 5 25
rect 3 -18 5 2
rect 3 -33 5 -28
<< polycontact >>
rect -1 -13 3 -9
<< metal1 >>
rect -9 28 17 33
rect -2 22 2 28
rect 6 -9 10 2
rect -7 -13 -1 -9
rect 6 -13 20 -9
rect 6 -18 10 -13
rect -2 -34 2 -28
rect -2 -38 10 -34
<< labels >>
rlabel metal1 -9 28 17 33 5 vdd
rlabel metal1 12 -11 20 -10 7 out
rlabel metal1 -6 -12 -4 -10 3 in
rlabel metal1 1 -37 6 -36 1 gnd
<< end >>
