* SPICE3 file created from dff_lbl.ext - technology: scmos

.include TSMC_180nm.txt
.option scale=0.09u
.global gnd Vdd

vdd vdd gnd 1.8

* Input Signals
Va2 d gnd PULSE(0 1.8 1.9ns 0ns 0ns 10ns 20ns)
VS clk gnd PULSE (0 1.8 2ns 0ns 0ns 3ns 6ns)

M1000 a_100_88# clk a_100_28# Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=240 ps=92
M1001 a_57_48# a_17_8# a_50_n12# w_44_38# CMOSP w=80 l=2
+  ad=480 pd=172 as=400 ps=170
M1002 dff_op a_100_88# vdd w_132_78# CMOSP w=40 l=2
+  ad=200 pd=90 as=1200 ps=520
M1003 a_17_48# d vdd w_4_38# CMOSP w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1004 a_57_n12# a_17_8# a_50_n12# Gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=200 ps=90
M1005 a_100_88# a_50_n12# vdd w_87_78# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1006 gnd clk a_57_n12# Gnd CMOSN w=40 l=2
+  ad=600 pd=280 as=0 ps=0
M1007 a_17_8# clk a_17_48# w_4_38# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1008 vdd clk a_57_48# w_44_38# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_100_28# a_50_n12# gnd Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 dff_op a_100_88# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1011 a_17_8# d gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 gnd a_50_n12# 0.05fF
C1 gnd a_100_88# 0.07fF
C2 vdd a_17_8# 0.09fF
C3 a_57_48# vdd 0.82fF
C4 w_132_78# dff_op 0.08fF
C5 a_17_48# w_4_38# 0.01fF
C6 vdd w_44_38# 0.42fF
C7 d clk 0.18fF
C8 a_50_n12# clk 0.49fF
C9 a_100_88# clk 0.08fF
C10 gnd a_100_28# 0.44fF
C11 d w_4_38# 0.14fF
C12 a_17_8# w_44_38# 0.14fF
C13 a_57_48# w_44_38# 0.01fF
C14 w_87_78# clk 0.36fF
C15 w_132_78# a_100_88# 0.09fF
C16 gnd a_17_8# 0.21fF
C17 dff_op a_100_88# 0.05fF
C18 vdd clk 0.02fF
C19 a_50_n12# a_57_n12# 0.44fF
C20 vdd w_4_38# 0.39fF
C21 w_132_78# vdd 0.19fF
C22 dff_op vdd 0.41fF
C23 a_17_8# clk 0.51fF
C24 clk w_44_38# 0.14fF
C25 vdd a_17_48# 0.82fF
C26 a_17_8# w_4_38# 0.25fF
C27 w_87_78# a_50_n12# 0.14fF
C28 w_87_78# a_100_88# 0.08fF
C29 vdd d 0.01fF
C30 a_17_48# a_17_8# 0.86fF
C31 vdd a_50_n12# 0.60fF
C32 a_100_88# vdd 0.41fF
C33 a_100_88# a_100_28# 0.41fF
C34 dff_op gnd 0.21fF
C35 w_87_78# vdd 0.30fF
C36 gnd a_57_n12# 0.44fF
C37 a_17_8# a_50_n12# 0.08fF
C38 a_57_48# a_50_n12# 0.82fF
C39 clk w_4_38# 0.14fF
C40 a_50_n12# w_44_38# 0.24fF
C41 a_57_n12# Gnd 0.01fF
C42 a_100_28# Gnd 0.01fF
C43 gnd Gnd 0.90fF
C44 dff_op Gnd 0.10fF
C45 a_100_88# Gnd 0.30fF
C46 vdd Gnd 0.32fF
C47 a_50_n12# Gnd 0.60fF
C48 a_17_8# Gnd 0.53fF
C49 clk Gnd 0.08fF
C50 d Gnd 0.08fF
C51 w_132_78# Gnd 1.51fF
C52 w_87_78# Gnd 1.62fF
C53 w_44_38# Gnd 3.38fF
C54 w_4_38# Gnd 3.28fF

.measure tran delay_dff_in
+TRIG v(clk) VAL=0.9 RISE=5
+TARG v(dff_op) VAL=0.9 FALL=2

.measure tran delay_dff_in_low_to_high
+TRIG v(clk) VAL=0.9 RISE=4
+TARG v(dff_op) VAL=0.9 RISE=2


.tran 1ps 50ns

.control
run
set color0 = white
set xbrushwidth = 3
set curplottitle = "Aditya_Peketi_2024122001_DFF"
plot v(dff_op) 2+v(d) 4+V(clk) 
.endc
