magic
tech scmos
timestamp 1731925082
<< nwell >>
rect 4 38 29 98
rect 42 39 67 99
rect 75 54 132 79
<< ntransistor >>
rect 15 8 17 28
rect 53 9 55 29
rect 84 21 104 23
<< ptransistor >>
rect 15 48 17 88
rect 53 49 55 89
rect 85 65 125 67
<< ndiffusion >>
rect 14 8 15 28
rect 17 8 18 28
rect 52 9 53 29
rect 55 9 56 29
rect 84 23 104 24
rect 84 20 104 21
<< pdiffusion >>
rect 14 48 15 88
rect 17 48 18 88
rect 52 49 53 89
rect 55 49 56 89
rect 85 67 125 68
rect 85 64 125 65
<< ndcontact >>
rect 10 8 14 28
rect 18 8 22 28
rect 48 9 52 29
rect 56 9 60 29
rect 84 24 104 28
rect 84 16 104 20
<< pdcontact >>
rect 10 48 14 88
rect 18 48 22 88
rect 48 49 52 89
rect 56 49 60 89
rect 85 68 125 72
rect 85 60 125 64
<< polysilicon >>
rect 15 88 17 106
rect 53 89 55 122
rect 78 65 85 67
rect 125 65 128 67
rect 15 28 17 48
rect 53 29 55 49
rect 77 21 84 23
rect 104 21 107 23
rect 15 5 17 8
rect 53 6 55 9
<< polycontact >>
rect 52 122 56 126
rect 14 106 18 110
rect 78 67 82 71
rect 77 17 81 21
<< metal1 >>
rect 56 122 142 126
rect 78 110 82 111
rect 18 106 82 110
rect 4 94 29 98
rect 44 97 48 106
rect 10 88 14 94
rect 44 93 52 97
rect 48 89 52 93
rect 78 71 82 106
rect 137 72 142 122
rect 125 68 142 72
rect 18 35 22 48
rect 56 38 60 49
rect 74 60 85 64
rect 74 39 78 60
rect 18 31 33 35
rect 18 28 22 31
rect 29 11 33 31
rect 56 34 73 38
rect 56 29 60 34
rect 10 4 14 8
rect 29 7 41 11
rect 4 0 29 4
rect 37 3 41 7
rect 74 28 78 32
rect 74 24 84 28
rect 137 20 142 68
rect 48 4 52 9
rect 77 4 81 17
rect 104 16 142 20
rect 48 3 81 4
rect 37 0 81 3
<< metal2 >>
rect 80 34 151 38
<< m123contact >>
rect 73 32 80 39
<< end >>
